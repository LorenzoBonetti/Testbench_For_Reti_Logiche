----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 12.12.2017 17:48:44
-- Design Name: 
-- Module Name: FSM_testbench - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
 
entity project_tb is
end project_tb;


architecture projecttb of project_tb is
constant c_CLOCK_PERIOD		: time := 15 ns;
signal   tb_done		: std_logic;
signal   mem_address		: std_logic_vector (15 downto 0) := (others => '0');
signal   tb_rst		    : std_logic := '0';
signal   tb_start		: std_logic := '0';
signal   tb_clk		    : std_logic := '0';
signal   mem_o_data,mem_i_data		: std_logic_vector (7 downto 0);
signal   enable_wire  		: std_logic;
signal   mem_we		: std_logic;

type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
--test # 1
signal RAM: ram_type := (2 => "00011000", 3 =>"00000111",4 => "00010101", 30 => "00000011", 31 => "00000011", 32 => "00000011", 33 => "00000011", 36 => "00000111", 37 => "00000111", 38 => "00000111", 39 => "00000111", 42 => "00001011", 43 => "00001011", 44 => "00001011", 45 => "00001011", 48 => "00001111", 54 => "00000011", 60 => "00000111", 66 => "00011111", 72 => "00011001", 78 => "00000011", 79 => "00000011", 80 => "00000011", 84 => "00000111", 85 => "00000111", 86 => "00000111", 90 => "00011111", 91 => "00011111", 92 => "00011111", 96 => "00011001", 102 => "00000011", 108 => "00000111", 114 => "00011111", 120 => "00011001", 126 => "00000011", 132 => "00000111", 133 => "00000111", 134 => "00000111", 135 => "00000111", 138 => "00001011", 139 => "00001011", 140 => "00001011", 141 => "00001011", 144 => "00001111", 145 => "00001111", 146 => "00001111", 147 => "00001111", others => (others =>'0'));
signal count : integer := 1;

component project_reti_logiche is 
    port (
            i_clk         : in  std_logic;
            i_start       : in  std_logic;
            i_rst         : in  std_logic;
            i_data       : in  std_logic_vector(7 downto 0); --1 byte
            o_address     : out std_logic_vector(15 downto 0); --16 bit addr: max size is 255*255 + 3 more for max x and y and thresh.
            o_done            : out std_logic;
            o_en         : out std_logic;
            o_we       : out std_logic;
            o_data            : out std_logic_vector (7 downto 0)
          );
end component project_reti_logiche;


begin 
	UUT: project_reti_logiche
	port map (
		  i_clk      	=> tb_clk,	
          i_start       => tb_start,
          i_rst      	=> tb_rst,
          i_data    	=> mem_o_data,
          o_address  	=> mem_address, 
          o_done      	=> tb_done,
          o_en   	=> enable_wire,
		  o_we 	=> mem_we,
          o_data    => mem_i_data
);

p_CLK_GEN : process is
  begin
    wait for c_CLOCK_PERIOD/2;
    tb_clk <= not tb_clk;
  end process p_CLK_GEN; 
  
  
MEM : process(tb_clk)
   begin
    if tb_clk'event and tb_clk = '1' then
    if enable_wire = '1' then
      if mem_we = '1' then
         RAM(conv_integer(mem_address))              <= mem_i_data;
         mem_o_data                      <= mem_i_data after 1 ns;
      else
        if tb_rst = '1' then
              if count = 1 then
              --test # 1
                RAM <= (2 => "00011000", 3 =>"00000111",4 => "00000000", 30 => "00000011", 31 => "00000011", 32 => "00000011", 33 => "00000011", 36 => "00000111", 37 => "00000111", 38 => "00000111", 39 => "00000111", 42 => "00001011", 43 => "00001011", 44 => "00001011", 45 => "00001011", 48 => "00001111", 54 => "00000011", 60 => "00000111", 66 => "00011111", 72 => "00011001", 78 => "00000011", 79 => "00000011", 80 => "00000011", 84 => "00000111", 85 => "00000111", 86 => "00000111", 90 => "00011111", 91 => "00011111", 92 => "00011111", 96 => "00011001", 102 => "00000011", 108 => "00000111", 114 => "00011111", 120 => "00011001", 126 => "00000011", 132 => "00000111", 133 => "00000111", 134 => "00000111", 135 => "00000111", 138 => "00001011", 139 => "00001011", 140 => "00001011", 141 => "00001011", 144 => "00001111", 145 => "00001111", 146 => "00001111", 147 => "00001111", others => (others =>'0'));
                count <= 2;
              elsif count = 2 then
              --test # 2
                RAM <= (2 => "00000000", 3 =>"00000111",4 => "00000000", 30 => "00000011", 31 => "00000011", 32 => "00000011", 33 => "00000011", 36 => "00000111", 37 => "00000111", 38 => "00000111", 39 => "00000111", 42 => "00001011", 43 => "00001011", 44 => "00001011", 45 => "00001011", 48 => "00001111", 54 => "00000011", 60 => "00000111", 66 => "00011111", 72 => "00011001", 78 => "00000011", 79 => "00000011", 80 => "00000011", 84 => "00000111", 85 => "00000111", 86 => "00000111", 90 => "00011111", 91 => "00011111", 92 => "00011111", 96 => "00011001", 102 => "00000011", 108 => "00000111", 114 => "00011111", 120 => "00011001", 126 => "00000011", 132 => "00000111", 133 => "00000111", 134 => "00000111", 135 => "00000111", 138 => "00001011", 139 => "00001011", 140 => "00001011", 141 => "00001011", 144 => "00001111", 145 => "00001111", 146 => "00001111", 147 => "00001111", others => (others =>'0'));
                count <= 3;
              elsif count = 3 then
              --test # 3
                RAM <= (2 => "00011000", 3 =>"00000000",4 => "00000000", 30 => "00000011", 31 => "00000011", 32 => "00000011", 33 => "00000011", 36 => "00000111", 37 => "00000111", 38 => "00000111", 39 => "00000111", 42 => "00001011", 43 => "00001011", 44 => "00001011", 45 => "00001011", 48 => "00001111", 54 => "00000011", 60 => "00000111", 66 => "00011111", 72 => "00011001", 78 => "00000011", 79 => "00000011", 80 => "00000011", 84 => "00000111", 85 => "00000111", 86 => "00000111", 90 => "00011111", 91 => "00011111", 92 => "00011111", 96 => "00011001", 102 => "00000011", 108 => "00000111", 114 => "00011111", 120 => "00011001", 126 => "00000011", 132 => "00000111", 133 => "00000111", 134 => "00000111", 135 => "00000111", 138 => "00001011", 139 => "00001011", 140 => "00001011", 141 => "00001011", 144 => "00001111", 145 => "00001111", 146 => "00001111", 147 => "00001111", others => (others =>'0'));
                count <= 4;  
              elsif count = 4 then
              --test # 4
                RAM <= (2 => "00000001", 3 =>"00000001",4 => "00100000",5 => "00010000",others => (others =>'0'));
                count <= 5;
            elsif count = 5 then
              --test # 5
                RAM <= (2 => "00000001", 3 =>"00000001",4 => "00010000",5 => "00010000",others => (others =>'0'));
                count <= 6;
            elsif count = 6 then
               --test # 6
                RAM <= (2 => "00000011", 3 =>"00000011",4 => "00010000",5 => "00010000",others => (others =>'0'));
                count <= 7;
            elsif count = 7 then 
               --test # 7
                RAM <= (2 => "00000011", 3 =>"00000011",4 => "00010000",13 => "00010000",others => (others =>'0'));
                mem_o_data <= "00000011" after 1 ns;
                count <= 8;
            elsif count = 8 then
               --test # 8
                RAM <= (2 => "00000110", 3 =>"00000100",4 => "00010000",11 => "00010000",12 => "00010000",15 => "00010000",16 => "00010000",others => (others =>'0'));
                mem_o_data <= "00000110" after 1 ns;
                count <= 9;
            elsif count = 9 then
               --test # 9
                RAM <= (2 => "00000110", 3 =>"00000100",4 => "00010000",6 => "00010000",12 => "00010000",24 => "00010000",others => (others =>'0'));
                count <= 10;
            elsif count = 10 then
               --test # 10
                RAM <= (2 => "11111111", 3 =>"11111111",4 => "00000000",others => (others =>'0'));
                count <= 11;
            elsif count = 11 then
               --test # 11
                RAM <= (2 => "11111111", 3 =>"11111111",4 => "11111111",others => (others =>'0'));
                count <= 12;
            elsif count = 12 then
               --test # 12
                RAM <= (2 => "00001101", 3 => "00001000", 4 => "00100001",  5 => "00000011", 6 => "00000010", 7 => "00000001", 8 => "00000000", 9 => "00000010", 10 => "00000010", 11 => "00000010", 12 => "00000000", 13 => "00000011", 14 => "00000010", 15 => "00000010", 16 => "00000010", 17 => "00000011", 18 => "00000010", 19 => "00000100", 20 => "00000111", 21 => "00000100", 22 => "00001011", 23 => "00001001", 24 => "00000011", 25 => "00001011", 26 => "00001100", 27 => "00000010", 28 => "00000110", 29 => "00000001", 30 => "00000111", 31 => "00000110", 32 => "00000101", 33 => "00001111", 34 => "00001001", 35 => "00001001", 36 => "00001101", 37 => "00000011", 38 => "00010000", 39 => "00011010", 40 => "00010110", 41 => "00011010", 42 => "00011011", 43 => "00100010", 44 => "00000110", 45 => "00001110", 46 => "00010010", 47 => "00000111", 48 => "00010011", 49 => "00000010", 50 => "00001111", 51 => "01111011", 52 => "00100111", 53 => "00010110", 54 => "00011100", 55 => "00001010", 56 => "00000000", 57 => "00000101", 58 => "00000011", 59 => "00000000", 60 => "00010001", 61 => "00011010", 62 => "00000001", 63 => "00010100", 64 => "00001010", 65 => "00101001", 66 => "00011001", 67 => "00011101", 68 => "00101001", 69 => "00010110", 70 => "00001010", 71 => "00000011", 72 => "00001101", 73 => "00010101", 74 => "00011011", 75 => "00110000", 76 => "00001111", 77 => "00000000", 78 => "00001010", 79 => "00010001", 80 => "00011001", 81 => "00001101", 82 => "01001011", 83 => "00000000", 84 => "00001111", 85 => "00010011", 86 => "00011101", 87 => "00010011", 88 => "00101101", 89 => "00000010", 90 => "00010100", 91 => "00010010", 92 => "00001001", 93 => "01001101", 94 => "01000000", 95 => "00011000", 96 => "00011110", 97 => "00010000", 98 => "00001101", 99 => "00001001", 100 => "00110100", 101 => "00000101", 102 => "00111111", 103 => "00000001", 104 => "00011111", 105 => "00111111", 106 => "00101101", 107 => "00010101", 108 => "00001001",others => (others =>'0'));
                count <= 13;
            elsif count =13  then
               --test # 13
                RAM <= (2 => "00001101", 3 => "00001000", 4 => "10110100",  5 => "00000011", 6 => "00000010", 7 => "00000001", 8 => "00000000", 9 => "00000010", 10 => "00000010", 11 => "00000010", 12 => "00000000", 13 => "00000011", 14 => "00000010", 15 => "00000010", 16 => "00000010", 17 => "00000011", 18 => "00000010", 19 => "00000100", 20 => "00000111", 21 => "00000100", 22 => "00001011", 23 => "00001001", 24 => "00000011", 25 => "00001011", 26 => "00001100", 27 => "00000010", 28 => "00000110", 29 => "00000001", 30 => "00000111", 31 => "00000110", 32 => "00000101", 33 => "00001111", 34 => "00001001", 35 => "00001001", 36 => "00001101", 37 => "00000011", 38 => "00010000", 39 => "00011010", 40 => "00010110", 41 => "00011010", 42 => "00011011", 43 => "00100010", 44 => "00000110", 45 => "00001110", 46 => "00010010", 47 => "00000111", 48 => "00010011", 49 => "00000010", 50 => "00001111", 51 => "01111011", 52 => "00100111", 53 => "00010110", 54 => "00011100", 55 => "00001010", 56 => "00000000", 57 => "00000101", 58 => "00000011", 59 => "00000000", 60 => "00010001", 61 => "00011010", 62 => "00000001", 63 => "00010100", 64 => "00001010", 65 => "00101001", 66 => "00011001", 67 => "00011101", 68 => "00101001", 69 => "00010110", 70 => "00001010", 71 => "00000011", 72 => "00001101", 73 => "00010101", 74 => "00011011", 75 => "00110000", 76 => "00001111", 77 => "00000000", 78 => "00001010", 79 => "00010001", 80 => "00011001", 81 => "00001101", 82 => "01001011", 83 => "00000000", 84 => "00001111", 85 => "00010011", 86 => "00011101", 87 => "00010011", 88 => "00101101", 89 => "00000010", 90 => "00010100", 91 => "00010010", 92 => "00001001", 93 => "01001101", 94 => "01000000", 95 => "00011000", 96 => "00011110", 97 => "00010000", 98 => "00001101", 99 => "00001001", 100 => "00110100", 101 => "00000101", 102 => "00111111", 103 => "00000001", 104 => "00011111", 105 => "00111111", 106 => "00101101", 107 => "00010101", 108 => "11001000", others => (others =>'0'));
                count <= 14;
            elsif count = 14  then
               --test # 14
                RAM <= (2 => "11111111", 3 =>"11111111",4 => "00000001", 30 => "00000011", 31 => "00000011", 32 => "00000011", 33 => "00000011", 36 => "00000111", 285 =>"00001000" , 291 =>"00001000" ,others => (others =>'0'));
                count <= 15;
            elsif count = 15 then
               --test # 15
                RAM <= (2 => "00001101", 3 => "00001000", 4 => "01100100",  5 => "00000011", 6 => "00000010", 7 => "00000001", 8 => "00000000", 9 => "11001000", 10 => "00000010", 11 => "00000010", 12 => "00000000", 13 => "00000011", 14 => "00000010", 15 => "00000010", 16 => "00000010", 17 => "00000011", 18 => "00000010", 19 => "00000100", 20 => "00000111", 21 => "00000100", 22 => "01110011", 23 => "00001001", 24 => "00000011", 25 => "00001011", 26 => "00001100", 27 => "00000010", 28 => "00000110", 29 => "00000001", 30 => "00000111", 31 => "00000110", 32 => "00000101", 33 => "00001111", 34 => "00001001", 35 => "10000100", 36 => "00001101", 37 => "00000011", 38 => "00010000", 39 => "00011010", 40 => "00010110", 41 => "00011010", 42 => "00011011", 43 => "00100010", 44 => "00000110", 45 => "00001110", 46 => "00010010", 47 => "00000111", 48 => "10111110", 49 => "00000010", 50 => "00001111", 51 => "00001100", 52 => "00100111", 53 => "00010110", 54 => "00011100", 55 => "00001010", 56 => "00000000", 57 => "00000101", 58 => "00000011", 59 => "00000000", 60 => "00010001", 61 => "11110111", 62 => "00000001", 63 => "00010100", 64 => "00001010", 65 => "00101001", 66 => "00011001", 67 => "00011101", 68 => "00101001", 69 => "00010110", 70 => "00001010", 71 => "00000011", 72 => "00001101", 73 => "00010101", 74 => "11011111", 75 => "00110000", 76 => "00001111", 77 => "00000000", 78 => "00001010", 79 => "00010001", 80 => "00011001", 81 => "00001101", 82 => "01001011", 83 => "00000000", 84 => "00001111", 85 => "00010011", 86 => "00011101", 87 => "10111110", 88 => "00101101", 89 => "00000010", 90 => "00010100", 91 => "00010010", 92 => "00001001", 93 => "01001101", 94 => "01000000", 95 => "00011000", 96 => "00011110", 97 => "00010000", 98 => "00001101", 99 => "00001001", 100 => "01111100", 101 => "00000101", 102 => "00111111", 103 => "00000001", 104 => "00011111", 105 => "00111111", 106 => "00101101", 107 => "00010101", 108 => "00001001", others => (others =>'0'));
                count <= 16;
            elsif count = 16 then
               --test # 16
                RAM <= (2 => "00001101", 3 => "00001000", 4 => "01101110",  5 => "00000011", 6 => "00000010", 7 => "00000001", 8 => "00000000", 9 => "00010100", 10 => "00000010", 11 => "00000010", 12 => "00000000", 13 => "00000011", 14 => "00000010", 15 => "00000010", 16 => "00000010", 17 => "00000011", 18 => "00000010", 19 => "00000100", 20 => "00000111", 21 => "00000100", 22 => "00001011", 23 => "00001001", 24 => "00000011", 25 => "00001011", 26 => "00001100", 27 => "00000010", 28 => "00000110", 29 => "00000001", 30 => "00000111", 31 => "00000110", 32 => "00000101", 33 => "00001111", 34 => "00001001", 35 => "10000100", 36 => "00001101", 37 => "00000011", 38 => "00010000", 39 => "00011010", 40 => "11011100", 41 => "00011010", 42 => "00011011", 43 => "00100010", 44 => "00000110", 45 => "00001110", 46 => "00010010", 47 => "00000111", 48 => "10111110", 49 => "00000010", 50 => "00001111", 51 => "00001100", 52 => "00100111", 53 => "00010110", 54 => "00011100", 55 => "00001010", 56 => "00000000", 57 => "00000101", 58 => "00000011", 59 => "00000000", 60 => "00010001", 61 => "11110111", 62 => "00000001", 63 => "00010100", 64 => "00001010", 65 => "00101001", 66 => "00011001", 67 => "00011101", 68 => "00101001", 69 => "00010110", 70 => "00001010", 71 => "00000011", 72 => "00001101", 73 => "00010101", 74 => "11011111", 75 => "00110000", 76 => "00001111", 77 => "00000000", 78 => "00001010", 79 => "00010001", 80 => "00011001", 81 => "00001101", 82 => "01001011", 83 => "00000000", 84 => "00001111", 85 => "00010011", 86 => "00011101", 87 => "00010011", 88 => "00101101", 89 => "00000010", 90 => "00010100", 91 => "00010010", 92 => "01111011", 93 => "01001101", 94 => "01000000", 95 => "00011000", 96 => "00011110", 97 => "00010000", 98 => "00001101", 99 => "00001001", 100 => "00000001", 101 => "00000101", 102 => "00111111", 103 => "00000001", 104 => "00011111", 105 => "00111111", 106 => "00101101", 107 => "00010101", 108 => "00001001", others => (others =>'0'));
                count <= 17;
            elsif count = 17 then
               --test # 17
                RAM <= (2 => "00001101", 3 => "00001000", 4 => "01111000",  5 => "00000011", 6 => "00000010", 7 => "00000001", 8 => "00000000", 9 => "00010100", 10 => "00000010", 11 => "00000010", 12 => "00000000", 13 => "00000011", 14 => "00000010", 15 => "00000010", 16 => "00000010", 17 => "01111001", 18 => "00000010", 19 => "00000100", 20 => "00000111", 21 => "00000100", 22 => "00001011", 23 => "00001001", 24 => "00000011", 25 => "00001011", 26 => "00001100", 27 => "00000010", 28 => "00000110", 29 => "00000001", 30 => "00000111", 31 => "00000110", 32 => "00000101", 33 => "10000010", 34 => "00001001", 35 => "10000100", 36 => "00001101", 37 => "00000011", 38 => "00010000", 39 => "00011010", 40 => "11011100", 41 => "00011010", 42 => "00011011", 43 => "00100010", 44 => "00000110", 45 => "00001110", 46 => "00010010", 47 => "00000111", 48 => "10111110", 49 => "00000010", 50 => "00001111", 51 => "00001100", 52 => "00100111", 53 => "00010110", 54 => "00011100", 55 => "00001010", 56 => "00000000", 57 => "00000101", 58 => "00000011", 59 => "00000000", 60 => "00010001", 61 => "11110111", 62 => "00000001", 63 => "00010100", 64 => "00001010", 65 => "00101001", 66 => "00011001", 67 => "00011101", 68 => "00101001", 69 => "00010110", 70 => "00001010", 71 => "00000011", 72 => "00001101", 73 => "00010101", 74 => "11011111", 75 => "00110000", 76 => "00001111", 77 => "00000000", 78 => "00001010", 79 => "00010001", 80 => "00011001", 81 => "00001101", 82 => "01001011", 83 => "00000000", 84 => "00001111", 85 => "00010011", 86 => "00011101", 87 => "00010011", 88 => "00101101", 89 => "00000010", 90 => "00010100", 91 => "00010010", 92 => "01111011", 93 => "01001101", 94 => "01000000", 95 => "00011000", 96 => "00011110", 97 => "00010000", 98 => "00001101", 99 => "00001001", 100 => "00000001", 101 => "00000101", 102 => "00111111", 103 => "00000001", 104 => "00011111", 105 => "00111111", 106 => "00101101", 107 => "00010101", 108 => "00001001", others => (others =>'0'));
                count <= 18;                  
            elsif count = 18 then
               --test # 18
                RAM <= (2 => "00001101", 3 => "00001000", 4 => "01111100",  5 => "00000011", 6 => "00000010", 7 => "00000001", 8 => "00000000", 9 => "00010100", 10 => "00000010", 11 => "00000010", 12 => "00000000", 13 => "00000011", 14 => "00000010", 15 => "00000010", 16 => "00000010", 17 => "00000001", 18 => "00000010", 19 => "00000100", 20 => "00000111", 21 => "00000100", 22 => "00001011", 23 => "00001001", 24 => "00000011", 25 => "00001011", 26 => "01111001", 27 => "00000010", 28 => "00000110", 29 => "00000001", 30 => "00000111", 31 => "00000110", 32 => "00000101", 33 => "10000010", 34 => "00001001", 35 => "10000100", 36 => "00001101", 37 => "00000011", 38 => "00010000", 39 => "00011010", 40 => "00010110", 41 => "00011010", 42 => "00011011", 43 => "00100010", 44 => "00000110", 45 => "00001110", 46 => "00010010", 47 => "00000111", 48 => "10111110", 49 => "00000010", 50 => "00001111", 51 => "00001100", 52 => "00100111", 53 => "00010110", 54 => "00011100", 55 => "00001010", 56 => "00000000", 57 => "00000101", 58 => "00000011", 59 => "00000000", 60 => "00010001", 61 => "11110111", 62 => "00000001", 63 => "00010100", 64 => "00001010", 65 => "00101001", 66 => "00011001", 67 => "00011101", 68 => "00101001", 69 => "00010110", 70 => "00001010", 71 => "00000011", 72 => "00001101", 73 => "00010101", 74 => "11011111", 75 => "00110000", 76 => "10011011", 77 => "00000000", 78 => "00001010", 79 => "00010001", 80 => "00011001", 81 => "00001101", 82 => "01001011", 83 => "00000000", 84 => "00001111", 85 => "00010011", 86 => "00011101", 87 => "00010011", 88 => "00101101", 89 => "00000010", 90 => "00010100", 91 => "00010010", 92 => "00001100", 93 => "01001101", 94 => "01000000", 95 => "00011000", 96 => "10000010", 97 => "00010000", 98 => "00001101", 99 => "10000110", 100 => "00000001", 101 => "00000101", 102 => "00111111", 103 => "00000001", 104 => "00011111", 105 => "00111111", 106 => "00101101", 107 => "00010101", 108 => "00001001", others => (others =>'0'));
                count <= 19;
            elsif count = 19 then
               --test # 19
                RAM <= (2 => "00001101", 3 => "00001000", 4 => "00101000",  5 => "00001101", 6 => "00000010", 7 => "00000001", 8 => "00000000", 9 => "00010100", 10 => "00000010", 11 => "00000010", 12 => "00000000", 13 => "00000011", 14 => "00000010", 15 => "00000010", 16 => "00000010", 17 => "00000001", 18 => "00000010", 19 => "00000100", 20 => "00000111", 21 => "00000100", 22 => "00001011", 23 => "00001001", 24 => "00000011", 25 => "00001011", 26 => "01111001", 27 => "00000010", 28 => "00000110", 29 => "00000001", 30 => "00000111", 31 => "00000110", 32 => "00000101", 33 => "10000010", 34 => "00001001", 35 => "10000100", 36 => "00001101", 37 => "00000011", 38 => "00010000", 39 => "00011010", 40 => "00010110", 41 => "00011010", 42 => "00011011", 43 => "00100010", 44 => "00000110", 45 => "00001110", 46 => "00010010", 47 => "00000111", 48 => "10111110", 49 => "00000010", 50 => "00001111", 51 => "00001100", 52 => "00100111", 53 => "00010110", 54 => "00011100", 55 => "00001010", 56 => "00000000", 57 => "00000101", 58 => "00000011", 59 => "00000000", 60 => "00010001", 61 => "11110111", 62 => "00000001", 63 => "00010100", 64 => "00001010", 65 => "00101001", 66 => "00011001", 67 => "00011101", 68 => "00101001", 69 => "00010110", 70 => "00001010", 71 => "00000011", 72 => "00001101", 73 => "00010101", 74 => "11011111", 75 => "00110000", 76 => "10011011", 77 => "00000000", 78 => "00001010", 79 => "00010001", 80 => "00011001", 81 => "00001101", 82 => "00000101", 83 => "00000000", 84 => "00001111", 85 => "00010011", 86 => "00011101", 87 => "00010011", 88 => "00101101", 89 => "00000010", 90 => "00010100", 91 => "00010010", 92 => "00001100", 93 => "01001101", 94 => "01000000", 95 => "00011000", 96 => "10000010", 97 => "00010000", 98 => "00001101", 99 => "10000110", 100 => "00000001", 101 => "00000101", 102 => "00111111", 103 => "00000001", 104 => "00011111", 105 => "00111111", 106 => "00101101", 107 => "00010101", 108 => "00001001", others => (others =>'0'));
                count <= 20;
            elsif count = 20 then
               --test # 20
                RAM <= (2 => "00010000", 3 => "00001011", 4 => "11001000",  5 => "00001101", 6 => "00000010", 7 => "00000001", 8 => "00000000", 9 => "00010100", 10 => "00000010", 11 => "00000010", 12 => "00000000", 13 => "00000011", 14 => "00000010", 15 => "00000010", 16 => "00000010", 17 => "00000001", 18 => "00000010", 19 => "00000001", 20 => "00000000", 21 => "00000010", 22 => "00000100", 23 => "00000111", 24 => "00000100", 25 => "00001011", 26 => "00001001", 27 => "00000011", 28 => "00001011", 29 => "01111001", 30 => "00000010", 31 => "00000110", 32 => "00000001", 33 => "00000111", 34 => "00000010", 35 => "00000001", 36 => "00000000", 37 => "00000110", 38 => "00000101", 39 => "10000010", 40 => "00001001", 41 => "10000100", 42 => "00001101", 43 => "00000011", 44 => "00010000", 45 => "00011010", 46 => "00010110", 47 => "00011010", 48 => "00011011", 49 => "00100010", 50 => "00000010", 51 => "00000001", 52 => "00000000", 53 => "00000110", 54 => "00001110", 55 => "00010010", 56 => "00000111", 57 => "10111110", 58 => "00000010", 59 => "00001111", 60 => "00001100", 61 => "00100111", 62 => "00010110", 63 => "00011100", 64 => "00001010", 65 => "00000000", 66 => "00000010", 67 => "00000001", 68 => "00000000", 69 => "00000101", 70 => "00000011", 71 => "00000000", 72 => "00010001", 73 => "11110111", 74 => "11101001", 75 => "00010100", 76 => "00001010", 77 => "00101001", 78 => "00011001", 79 => "00011101", 80 => "00101001", 81 => "00010110", 82 => "00000010", 83 => "00000001", 84 => "00000000", 85 => "00001010", 86 => "00000011", 87 => "00001101", 88 => "00010101", 89 => "11011111", 90 => "11100111", 91 => "10011011", 92 => "00000000", 93 => "00001010", 94 => "00010001", 95 => "00011001", 96 => "00001101", 97 => "00000101", 98 => "00000010", 99 => "00000001", 100 => "00000000", 101 => "00000000", 102 => "00001111", 103 => "00010011", 104 => "00011101", 105 => "00010011", 106 => "00101101", 107 => "00000010", 108 => "00010100", 109 => "00010010", 110 => "00001100", 111 => "01001101", 112 => "01000000", 113 => "00011000", 114 => "00000010", 115 => "00000001", 116 => "00000000", 117 => "00000000", 118 => "00001111", 119 => "00010011", 120 => "00011101", 121 => "00010011", 122 => "00101101", 123 => "00000010", 124 => "00010100", 125 => "00010010", 126 => "00001100", 127 => "01001101", 128 => "01000000", 129 => "00011000", 130 => "00000010", 131 => "00000001", 132 => "00000000", 133 => "00000000", 134 => "00001111", 135 => "00010011", 136 => "00011101", 137 => "00010011", 138 => "00101101", 139 => "00000010", 140 => "00010100", 141 => "00010010", 142 => "00001100", 143 => "01001101", 144 => "01000000", 145 => "00011000", 146 => "00000010", 147 => "00000001", 148 => "00000000", 149 => "00000000", 150 => "00001111", 151 => "00010011", 152 => "00011101", 153 => "00010011", 154 => "00101101", 155 => "00000010", 156 => "00010100", 157 => "00010010", 158 => "00001100", 159 => "01001101", 160 => "01000000", 161 => "00011000", 162 => "00000010", 163 => "00000001", 164 => "00000000", 165 => "10000010", 166 => "00010000", 167 => "00001101", 168 => "10000110", 169 => "00000001", 170 => "00000101", 171 => "00111111", 172 => "00000001", 173 => "00011111", 174 => "00111111", 175 => "00101101", 176 => "00010101", 177 => "00001001", 178 => "00000010", 179 => "00000001", 180 => "00000000", others => (others =>'0'));
                count <= 21;
            elsif count = 21 then
               --test # 21
                RAM <= (2 => "00010000", 3 => "00001011", 4 => "00001010",  5 => "00001101", 6 => "00000010", 7 => "00000001", 8 => "00000000", 9 => "00010100", 10 => "00000010", 11 => "00000010", 12 => "00000000", 13 => "00000011", 14 => "01111011", 15 => "00000010", 16 => "00000010", 17 => "00000001", 18 => "11011110", 19 => "00000001", 20 => "00000000", 21 => "00000010", 22 => "00000100", 23 => "00000111", 24 => "00000100", 25 => "00001011", 26 => "00001001", 27 => "00000011", 28 => "00001011", 29 => "01111001", 30 => "00000010", 31 => "00000110", 32 => "00000001", 33 => "00000111", 34 => "00000010", 35 => "00000001", 36 => "00000000", 37 => "00000110", 38 => "00000101", 39 => "10000010", 40 => "00001001", 41 => "10000100", 42 => "00001101", 43 => "00000011", 44 => "00010000", 45 => "00011010", 46 => "00010110", 47 => "00011010", 48 => "00011011", 49 => "00100010", 50 => "00000010", 51 => "00000011", 52 => "00000000", 53 => "00000110", 54 => "00001100", 55 => "00010010", 56 => "00000111", 57 => "10111110", 58 => "00000010", 59 => "00001111", 60 => "00001100", 61 => "00100111", 62 => "00010110", 63 => "00011100", 64 => "00001010", 65 => "00000000", 66 => "00000010", 67 => "00000001", 68 => "00000000", 69 => "00000101", 70 => "00011110", 71 => "00000000", 72 => "00010001", 73 => "11110111", 74 => "00010111", 75 => "00010100", 76 => "00001010", 77 => "00101001", 78 => "00011001", 79 => "00011101", 80 => "00101001", 81 => "00010110", 82 => "00000010", 83 => "00000001", 84 => "00000000", 85 => "00001010", 86 => "00001100", 87 => "00001101", 88 => "00010101", 89 => "00010110", 90 => "11100111", 91 => "10011011", 92 => "00000000", 93 => "00001010", 94 => "00010001", 95 => "00011001", 96 => "00001101", 97 => "00110010", 98 => "00000010", 99 => "00000001", 100 => "00000100", 101 => "00000000", 102 => "00001111", 103 => "00010011", 104 => "00011101", 105 => "00010011", 106 => "00101101", 107 => "00000010", 108 => "00010100", 109 => "00010010", 110 => "00001100", 111 => "01001101", 112 => "01000000", 113 => "00011000", 114 => "00000010", 115 => "00000011", 116 => "00000000", 117 => "00000000", 118 => "00001111", 119 => "00010011", 120 => "00011101", 121 => "00010011", 122 => "00101101", 123 => "00000010", 124 => "00010100", 125 => "00100010", 126 => "00001100", 127 => "01001101", 128 => "01000000", 129 => "00011000", 130 => "00000010", 131 => "00000001", 132 => "00000000", 133 => "00000000", 134 => "00001111", 135 => "00010011", 136 => "00011101", 137 => "00010011", 138 => "00101101", 139 => "00000010", 140 => "00010100", 141 => "00010010", 142 => "00001100", 143 => "01001101", 144 => "01000000", 145 => "00011000", 146 => "00000010", 147 => "00000001", 148 => "00000110", 149 => "00000000", 150 => "00001111", 151 => "00010011", 152 => "00011101", 153 => "00010011", 154 => "00101101", 155 => "00000010", 156 => "00010100", 157 => "00010010", 158 => "00001100", 159 => "01001101", 160 => "01000000", 161 => "00011000", 162 => "00000010", 163 => "00001100", 164 => "00000000", 165 => "10000010", 166 => "00010000", 167 => "00001101", 168 => "10000110", 169 => "00000001", 170 => "00000101", 171 => "00111111", 172 => "00000001", 173 => "00011111", 174 => "00111111", 175 => "00101101", 176 => "00010101", 177 => "00001001", 178 => "00000010", 179 => "00000001", 180 => "00000000", others => (others =>'0'));
                count <= 22;
            elsif count = 22 then
               --test # 22
                RAM <= (2 => "00010000", 3 => "00001011", 4 => "01111100",  5 => "00001101", 6 => "00000010", 7 => "00000001", 8 => "00000000", 9 => "00010100", 10 => "00000010", 11 => "00000010", 12 => "00000000", 13 => "00000011", 14 => "00001100", 15 => "00000010", 16 => "00000010", 17 => "00000001", 18 => "00010110", 19 => "00000001", 20 => "00000000", 21 => "00000010", 22 => "00000100", 23 => "00000111", 24 => "00000100", 25 => "00001011", 26 => "00001001", 27 => "00000011", 28 => "00001011", 29 => "01111001", 30 => "00000010", 31 => "00000110", 32 => "00000001", 33 => "00000111", 34 => "00000010", 35 => "00000001", 36 => "00000000", 37 => "00000110", 38 => "00000101", 39 => "10000010", 40 => "00001001", 41 => "10000100", 42 => "00001101", 43 => "00000011", 44 => "00010000", 45 => "00011010", 46 => "00010110", 47 => "00011010", 48 => "00011011", 49 => "00100010", 50 => "00000010", 51 => "00000011", 52 => "00000000", 53 => "00000110", 54 => "00001100", 55 => "00010010", 56 => "00000111", 57 => "10111110", 58 => "00000010", 59 => "00001111", 60 => "00001100", 61 => "00100111", 62 => "00010110", 63 => "00011100", 64 => "00001010", 65 => "00000000", 66 => "00000010", 67 => "00000001", 68 => "00000000", 69 => "00000101", 70 => "00011110", 71 => "00000000", 72 => "00010001", 73 => "11110111", 74 => "00010111", 75 => "00010100", 76 => "00001010", 77 => "00101001", 78 => "00011001", 79 => "00011101", 80 => "00101001", 81 => "00010110", 82 => "00000010", 83 => "00000001", 84 => "00000000", 85 => "00001010", 86 => "00001100", 87 => "00001101", 88 => "00010101", 89 => "00010110", 90 => "11100111", 91 => "10011011", 92 => "00000000", 93 => "00001010", 94 => "00010001", 95 => "00011001", 96 => "00001101", 97 => "00110010", 98 => "00000010", 99 => "00000001", 100 => "00000100", 101 => "00000000", 102 => "00001111", 103 => "00010011", 104 => "00011101", 105 => "00010011", 106 => "00101101", 107 => "00000010", 108 => "00010100", 109 => "00010010", 110 => "00001100", 111 => "01001101", 112 => "01000000", 113 => "00011000", 114 => "00000010", 115 => "00000011", 116 => "00000000", 117 => "00000000", 118 => "00001111", 119 => "00010011", 120 => "00011101", 121 => "00010011", 122 => "00101101", 123 => "00000010", 124 => "00010100", 125 => "00100010", 126 => "00001100", 127 => "01001101", 128 => "01000000", 129 => "00011000", 130 => "00000010", 131 => "00000001", 132 => "00000000", 133 => "00000000", 134 => "00001111", 135 => "00010011", 136 => "00011101", 137 => "00010011", 138 => "00101101", 139 => "00000010", 140 => "00010100", 141 => "00010010", 142 => "00001100", 143 => "01001101", 144 => "01000000", 145 => "00011000", 146 => "00000010", 147 => "00000001", 148 => "00000110", 149 => "00000000", 150 => "00001111", 151 => "00010011", 152 => "00011101", 153 => "00010011", 154 => "00101101", 155 => "00000010", 156 => "00010100", 157 => "00010010", 158 => "00001100", 159 => "01001101", 160 => "01000000", 161 => "00011000", 162 => "00000010", 163 => "00001100", 164 => "00000000", 165 => "00001101", 166 => "00010000", 167 => "00001101", 168 => "10000110", 169 => "00000001", 170 => "00000101", 171 => "00111111", 172 => "00000001", 173 => "00011111", 174 => "00111111", 175 => "00101101", 176 => "00010101", 177 => "00001001", 178 => "00000010", 179 => "00000001", 180 => "00000000", others => (others =>'0'));
                count <= 23;
            elsif count = 23 then
               --test # 23
                RAM <= (2 => "00010000", 3 => "00001011", 4 => "11111010",  5 => "00001101", 6 => "00000010", 7 => "00000001", 8 => "00000000", 9 => "00010100", 10 => "00000010", 11 => "00000010", 12 => "00000000", 13 => "00000011", 14 => "00001100", 15 => "00000010", 16 => "00000010", 17 => "00000001", 18 => "00010110", 19 => "00000001", 20 => "00000000", 21 => "00000010", 22 => "00000100", 23 => "00000111", 24 => "00000100", 25 => "00001011", 26 => "00001001", 27 => "00000011", 28 => "00001011", 29 => "01111001", 30 => "00000010", 31 => "00000110", 32 => "00000001", 33 => "00000111", 34 => "00000010", 35 => "00000001", 36 => "00000000", 37 => "00000110", 38 => "00000101", 39 => "10000010", 40 => "00001001", 41 => "10000100", 42 => "00001101", 43 => "00000011", 44 => "00010000", 45 => "00011010", 46 => "00010110", 47 => "00011010", 48 => "00011011", 49 => "00100010", 50 => "00000010", 51 => "00000011", 52 => "00000000", 53 => "00000110", 54 => "00001100", 55 => "00010010", 56 => "00000111", 57 => "10111110", 58 => "00000010", 59 => "00001111", 60 => "00001100", 61 => "00100111", 62 => "00010110", 63 => "00011100", 64 => "00001010", 65 => "00000000", 66 => "00000010", 67 => "00000001", 68 => "00000000", 69 => "00000101", 70 => "00011110", 71 => "00000000", 72 => "00010001", 73 => "11110111", 74 => "00010111", 75 => "00010100", 76 => "00001010", 77 => "00101001", 78 => "00011001", 79 => "00011101", 80 => "00101001", 81 => "00010110", 82 => "00000010", 83 => "00000001", 84 => "00000000", 85 => "00001010", 86 => "00001100", 87 => "00001101", 88 => "00010101", 89 => "00010110", 90 => "11100111", 91 => "10011011", 92 => "00000000", 93 => "00001010", 94 => "00010001", 95 => "00011001", 96 => "00001101", 97 => "00110010", 98 => "00000010", 99 => "00000001", 100 => "00000100", 101 => "00000000", 102 => "00001111", 103 => "00010011", 104 => "00011101", 105 => "00010011", 106 => "00101101", 107 => "00000010", 108 => "00010100", 109 => "00010010", 110 => "00001100", 111 => "01001101", 112 => "01000000", 113 => "00011000", 114 => "00000010", 115 => "00000011", 116 => "00000000", 117 => "00000000", 118 => "00001111", 119 => "00010011", 120 => "00011101", 121 => "00010011", 122 => "00101101", 123 => "00000010", 124 => "00010100", 125 => "00100010", 126 => "00001100", 127 => "01001101", 128 => "01000000", 129 => "00011000", 130 => "00000010", 131 => "00000001", 132 => "00000000", 133 => "00000000", 134 => "00001111", 135 => "00010011", 136 => "00011101", 137 => "00010011", 138 => "00101101", 139 => "00000010", 140 => "00010100", 141 => "00010010", 142 => "00001100", 143 => "01001101", 144 => "01000000", 145 => "00011000", 146 => "00000010", 147 => "00000001", 148 => "00000110", 149 => "00000000", 150 => "00001111", 151 => "00010011", 152 => "00011101", 153 => "00010011", 154 => "00101101", 155 => "00000010", 156 => "00010100", 157 => "00010010", 158 => "00001100", 159 => "01001101", 160 => "01000000", 161 => "00011000", 162 => "00000010", 163 => "00001100", 164 => "00000000", 165 => "00001101", 166 => "00010000", 167 => "00001101", 168 => "10000110", 169 => "00000001", 170 => "00000101", 171 => "00111111", 172 => "00000001", 173 => "00011111", 174 => "00111111", 175 => "00101101", 176 => "00010101", 177 => "00001001", 178 => "00000010", 179 => "00000001", 180 => "00000000", others => (others =>'0'));
                count <= 24;
            elsif count = 24 then
               --test # 24
                RAM <= (2 => "00010000", 3 => "00001011", 4 => "11111010",  5 => "00001101", 6 => "00000010", 7 => "00000001", 8 => "00000000", 9 => "00010100", 10 => "00000010", 11 => "00000010", 12 => "00000000", 13 => "00000011", 14 => "00001100", 15 => "00000010", 16 => "00000010", 17 => "00000001", 18 => "00010110", 19 => "00000001", 20 => "00000000", 21 => "00000010", 22 => "00000100", 23 => "00000111", 24 => "00000100", 25 => "00001011", 26 => "00001001", 27 => "00000011", 28 => "00001011", 29 => "01111001", 30 => "00000010", 31 => "00000110", 32 => "00000001", 33 => "00000111", 34 => "00000010", 35 => "00000001", 36 => "00000000", 37 => "00000110", 38 => "00000101", 39 => "10000010", 40 => "00001001", 41 => "10000100", 42 => "00001101", 43 => "00000011", 44 => "00010000", 45 => "00011010", 46 => "00010110", 47 => "00011010", 48 => "00011011", 49 => "00100010", 50 => "00000010", 51 => "00000011", 52 => "00000000", 53 => "00000110", 54 => "00001100", 55 => "00010010", 56 => "00000111", 57 => "10111110", 58 => "00000010", 59 => "00001111", 60 => "00001100", 61 => "00100111", 62 => "00010110", 63 => "00011100", 64 => "00001010", 65 => "00000000", 66 => "00000010", 67 => "00000001", 68 => "00000000", 69 => "00000101", 70 => "00011110", 71 => "00000000", 72 => "00010001", 73 => "11110111", 74 => "00010111", 75 => "00010100", 76 => "00001010", 77 => "00101001", 78 => "00011001", 79 => "00011101", 80 => "00101001", 81 => "00010110", 82 => "00000010", 83 => "00000001", 84 => "00000000", 85 => "11111010", 86 => "11111010", 87 => "11111010", 88 => "11111010", 89 => "11111010", 90 => "11111010", 91 => "11111010", 92 => "11111010", 93 => "11111010", 94 => "11111010", 95 => "11111010", 96 => "11111010", 97 => "11111010", 98 => "11111010", 99 => "11111010", 100 => "11111010", 101 => "00000000", 102 => "00001111", 103 => "00010011", 104 => "00011101", 105 => "00010011", 106 => "00101101", 107 => "00000010", 108 => "00010100", 109 => "00010010", 110 => "00001100", 111 => "01001101", 112 => "01000000", 113 => "00011000", 114 => "00000010", 115 => "00000011", 116 => "00000000", 117 => "00000000", 118 => "00001111", 119 => "00010011", 120 => "00011101", 121 => "00010011", 122 => "00101101", 123 => "00000010", 124 => "00010100", 125 => "00100010", 126 => "00001100", 127 => "01001101", 128 => "01000000", 129 => "00011000", 130 => "00000010", 131 => "00000001", 132 => "00000000", 133 => "00000000", 134 => "00001111", 135 => "00010011", 136 => "00011101", 137 => "00010011", 138 => "00101101", 139 => "00000010", 140 => "00010100", 141 => "00010010", 142 => "00001100", 143 => "01001101", 144 => "01000000", 145 => "00011000", 146 => "00000010", 147 => "00000001", 148 => "00000110", 149 => "00000000", 150 => "00001111", 151 => "00010011", 152 => "00011101", 153 => "00010011", 154 => "00101101", 155 => "00000010", 156 => "00010100", 157 => "00010010", 158 => "00001100", 159 => "01001101", 160 => "01000000", 161 => "00011000", 162 => "00000010", 163 => "00001100", 164 => "00000000", 165 => "00001101", 166 => "00010000", 167 => "00001101", 168 => "10000110", 169 => "00000001", 170 => "00000101", 171 => "00111111", 172 => "00000001", 173 => "00011111", 174 => "00111111", 175 => "00101101", 176 => "00010101", 177 => "00001001", 178 => "00000010", 179 => "00000001", 180 => "00000000", others => (others =>'0'));
                count <= 25;
            elsif count = 25 then
               --test # 25
                RAM <= (2 => "00010000", 3 => "00001011", 4 => "11110111",  5 => "00001101", 6 => "00000010", 7 => "00000001", 8 => "00000000", 9 => "00010100", 10 => "00000010", 11 => "00000010", 12 => "00000000", 13 => "00000011", 14 => "00001100", 15 => "00000010", 16 => "00000010", 17 => "00000001", 18 => "00010110", 19 => "00000001", 20 => "00000000", 21 => "00000010", 22 => "00000100", 23 => "00000111", 24 => "00000100", 25 => "00001011", 26 => "00001001", 27 => "00000011", 28 => "00001011", 29 => "01111001", 30 => "00000010", 31 => "00000110", 32 => "00000001", 33 => "00000111", 34 => "00000010", 35 => "00000001", 36 => "00000000", 37 => "00000110", 38 => "00000101", 39 => "10000010", 40 => "00001001", 41 => "10000100", 42 => "00001101", 43 => "00000011", 44 => "00010000", 45 => "00011010", 46 => "00010110", 47 => "00011010", 48 => "00011011", 49 => "00100010", 50 => "00000010", 51 => "00000011", 52 => "00000000", 53 => "00000110", 54 => "00001100", 55 => "00010010", 56 => "00000111", 57 => "10111110", 58 => "00000010", 59 => "00001111", 60 => "00001100", 61 => "00100111", 62 => "00010110", 63 => "00011100", 64 => "00001010", 65 => "00000000", 66 => "00000010", 67 => "00000001", 68 => "00000000", 69 => "00000101", 70 => "00011110", 71 => "00000000", 72 => "00010001", 73 => "11110111", 74 => "00010111", 75 => "00010100", 76 => "00001010", 77 => "00101001", 78 => "00011001", 79 => "00011101", 80 => "00101001", 81 => "00010110", 82 => "00000010", 83 => "00000001", 84 => "00000000", 85 => "00000101", 86 => "00011110", 87 => "00000000", 88 => "00010001", 89 => "11110111", 90 => "00010111", 91 => "00010100", 92 => "00001010", 93 => "00101001", 94 => "00011001", 95 => "00011101", 96 => "00101001", 97 => "00010110", 98 => "00000010", 99 => "00000001", 100 => "00000000", 101 => "00000000", 102 => "00001111", 103 => "00010011", 104 => "00011101", 105 => "00010011", 106 => "00101101", 107 => "00000010", 108 => "00010100", 109 => "00010010", 110 => "00001100", 111 => "01001101", 112 => "01000000", 113 => "00011000", 114 => "00000010", 115 => "00000011", 116 => "00000000", 117 => "00000000", 118 => "00001111", 119 => "00010011", 120 => "00011101", 121 => "00010011", 122 => "00101101", 123 => "00000010", 124 => "00010100", 125 => "00100010", 126 => "00001100", 127 => "01001101", 128 => "01000000", 129 => "00011000", 130 => "00000010", 131 => "00000001", 132 => "00000000", 133 => "00000000", 134 => "00001111", 135 => "00010011", 136 => "00011101", 137 => "00010011", 138 => "00101101", 139 => "00000010", 140 => "00010100", 141 => "00010010", 142 => "00001100", 143 => "01001101", 144 => "01000000", 145 => "00011000", 146 => "00000010", 147 => "00000001", 148 => "00000110", 149 => "00000000", 150 => "00001111", 151 => "00010011", 152 => "00011101", 153 => "00010011", 154 => "00101101", 155 => "00000010", 156 => "00010100", 157 => "00010010", 158 => "00001100", 159 => "01001101", 160 => "01000000", 161 => "00011000", 162 => "00000010", 163 => "00001100", 164 => "00000000", 165 => "00001101", 166 => "00010000", 167 => "00001101", 168 => "10000110", 169 => "00000001", 170 => "00000101", 171 => "00111111", 172 => "00000001", 173 => "00011111", 174 => "00111111", 175 => "00101101", 176 => "00010101", 177 => "00001001", 178 => "00000010", 179 => "00000001", 180 => "00000000", others => (others =>'0'));
                count <= 26;
            elsif count = 26 then
               --test # 26
                RAM <= (2 => "00010100", 3 => "00001110", 4 => "00001101",  5 => "00000001", 6 => "00010110", 7 => "00000001", 8 => "00000000", 9 => "00010100", 10 => "00000010", 11 => "00000010", 12 => "00000000", 13 => "00000011", 14 => "00001100", 15 => "00000010", 16 => "00000010", 17 => "00000001", 18 => "00010110", 19 => "00000001", 20 => "00000110", 21 => "01001101", 22 => "01000000", 23 => "00011000", 24 => "00000010", 25 => "00000010", 26 => "00000100", 27 => "00000111", 28 => "00000100", 29 => "00001011", 30 => "00001001", 31 => "00000011", 32 => "00001011", 33 => "01111001", 34 => "00000010", 35 => "00000110", 36 => "00000001", 37 => "00000111", 38 => "00000010", 39 => "00000001", 40 => "00000000", 41 => "00000011", 42 => "00010000", 43 => "00011010", 44 => "00010110", 45 => "00000110", 46 => "00000101", 47 => "10000010", 48 => "00001001", 49 => "10000100", 50 => "00001101", 51 => "00000011", 52 => "00010000", 53 => "00011010", 54 => "00010110", 55 => "00011010", 56 => "00011011", 57 => "00100010", 58 => "00000010", 59 => "00000011", 60 => "00000011", 61 => "01001101", 62 => "01000000", 63 => "00011000", 64 => "00000010", 65 => "00000110", 66 => "00001100", 67 => "00010010", 68 => "00000111", 69 => "10111110", 70 => "00000010", 71 => "00001111", 72 => "00001100", 73 => "00100111", 74 => "00010110", 75 => "00011100", 76 => "00001010", 77 => "00000000", 78 => "00000010", 79 => "00000001", 80 => "00000000", 81 => "00010011", 82 => "00101101", 83 => "00000010", 84 => "00010100", 85 => "00000101", 86 => "00011110", 87 => "00000000", 88 => "00010001", 89 => "11110111", 90 => "00010111", 91 => "00010100", 92 => "00001010", 93 => "00101001", 94 => "01000010", 95 => "00011101", 96 => "00101001", 97 => "00010110", 98 => "00000010", 99 => "00000001", 100 => "00000001", 101 => "00000011", 102 => "00010000", 103 => "00011010", 104 => "00010110", 105 => "00000101", 106 => "00011110", 107 => "00000000", 108 => "00010001", 109 => "11110111", 110 => "00010111", 111 => "00010100", 112 => "00001010", 113 => "00101001", 114 => "00011001", 115 => "00011101", 116 => "00101001", 117 => "00010110", 118 => "00000010", 119 => "00000001", 120 => "00000000", 121 => "01001101", 122 => "01000000", 123 => "00011000", 124 => "00000010", 125 => "00000000", 126 => "00001111", 127 => "00010011", 128 => "00011101", 129 => "00010011", 130 => "00101101", 131 => "00000010", 132 => "00000001", 133 => "00010010", 134 => "00001100", 135 => "01001101", 136 => "01000000", 137 => "00011000", 138 => "00000010", 139 => "00000011", 140 => "00000000", 141 => "00000011", 142 => "00010000", 143 => "00011010", 144 => "00010110", 145 => "00000010", 146 => "00000100", 147 => "00000111", 148 => "00000100", 149 => "00001011", 150 => "00001001", 151 => "00000011", 152 => "00001011", 153 => "01111001", 154 => "00000010", 155 => "00000110", 156 => "00000001", 157 => "00000111", 158 => "00000010", 159 => "00000001", 160 => "00000000", 161 => "00000011", 162 => "00010000", 163 => "00011010", 164 => "00010110", 165 => "00000101", 166 => "00011110", 167 => "00000000", 168 => "00010001", 169 => "11110111", 170 => "00010111", 171 => "00010100", 172 => "00001010", 173 => "00101001", 174 => "00011001", 175 => "00011101", 176 => "00101001", 177 => "00010110", 178 => "00000010", 179 => "00000001", 180 => "00000010", 181 => "01001101", 182 => "01000000", 183 => "00011000", 184 => "00000010", 185 => "00000000", 186 => "00001111", 187 => "00010011", 188 => "00011101", 189 => "00010011", 190 => "00101101", 191 => "00000010", 192 => "00010100", 193 => "00010010", 194 => "00001100", 195 => "00001100", 196 => "01000000", 197 => "00011000", 198 => "00000010", 199 => "00001100", 200 => "00000000", 201 => "00000011", 202 => "00010000", 203 => "00011010", 204 => "00010110", 205 => "00000000", 206 => "00001111", 207 => "00010011", 208 => "00011101", 209 => "00010011", 210 => "00101101", 211 => "00000010", 212 => "00010110", 213 => "00100010", 214 => "00001100", 215 => "00101011", 216 => "01000000", 217 => "00011000", 218 => "00000010", 219 => "00000001", 220 => "00000000", 221 => "00000011", 222 => "00010000", 223 => "00011010", 224 => "00010110", 225 => "00000000", 226 => "00001111", 227 => "00010011", 228 => "00011101", 229 => "00010011", 230 => "00101101", 231 => "00000010", 232 => "00010100", 233 => "00010010", 234 => "00001100", 235 => "01001101", 236 => "01000000", 237 => "00011000", 238 => "00000010", 239 => "00000001", 240 => "00000110", 241 => "00010011", 242 => "00101101", 243 => "00000010", 244 => "00010100", 245 => "00000001", 246 => "00001111", 247 => "00010011", 248 => "00011101", 249 => "00010011", 250 => "00101101", 251 => "00000010", 252 => "00010100", 253 => "00010010", 254 => "00001100", 255 => "00001100", 256 => "01000000", 257 => "00011000", 258 => "00000010", 259 => "00001100", 260 => "00000000", 261 => "00000011", 262 => "00010000", 263 => "00011010", 264 => "00010110", 265 => "00000001", 266 => "00001111", 267 => "00001101", 268 => "00000001", 269 => "00000001", 270 => "00000101", 271 => "00000011", 272 => "00000001", 273 => "00000001", 274 => "00000011", 275 => "00000101", 276 => "00000001", 277 => "00001001", 278 => "00000010", 279 => "00000001", 280 => "00000100", 281 => "00000011", 282 => "00000110", 283 => "00000110", 284 => "00010110", others => (others =>'0'));
                count <= 27;
            elsif count = 27 then
               --test # 27
                RAM <= (2 => "00010100", 3 => "00001110", 4 => "11011110",  5 => "00000001", 6 => "00010110", 7 => "00000001", 8 => "00000000", 9 => "00010100", 10 => "00000010", 11 => "00000010", 12 => "00000000", 13 => "00000011", 14 => "00001100", 15 => "00000010", 16 => "00000010", 17 => "00000001", 18 => "00010110", 19 => "00000001", 20 => "00000110", 21 => "01001101", 22 => "01000000", 23 => "11110000", 24 => "00000010", 25 => "11011111", 26 => "00000100", 27 => "00000111", 28 => "00000100", 29 => "00001011", 30 => "00001001", 31 => "00000011", 32 => "00001011", 33 => "01111001", 34 => "00000010", 35 => "00000110", 36 => "00000001", 37 => "00000111", 38 => "00000010", 39 => "00000001", 40 => "00000000", 41 => "00000011", 42 => "00010000", 43 => "00011010", 44 => "00010110", 45 => "00000110", 46 => "00000101", 47 => "10000010", 48 => "00001001", 49 => "10000100", 50 => "00001101", 51 => "00000011", 52 => "00010000", 53 => "00011010", 54 => "00010110", 55 => "00011010", 56 => "00011011", 57 => "00100010", 58 => "00000010", 59 => "00000011", 60 => "00000011", 61 => "01001101", 62 => "01000000", 63 => "00011000", 64 => "00000010", 65 => "00000110", 66 => "00001100", 67 => "00010010", 68 => "00000111", 69 => "10111110", 70 => "00000010", 71 => "00001111", 72 => "00001100", 73 => "00100111", 74 => "00010110", 75 => "00011100", 76 => "00001010", 77 => "00000000", 78 => "00000010", 79 => "00000001", 80 => "00000000", 81 => "00010011", 82 => "00101101", 83 => "00000010", 84 => "00010100", 85 => "00000101", 86 => "00011110", 87 => "00000000", 88 => "00010001", 89 => "11110111", 90 => "00010111", 91 => "00010100", 92 => "00001010", 93 => "00101001", 94 => "01000010", 95 => "00011101", 96 => "00101001", 97 => "00010110", 98 => "00000010", 99 => "00000001", 100 => "00000001", 101 => "00000011", 102 => "00010000", 103 => "00011010", 104 => "00010110", 105 => "00000101", 106 => "00011110", 107 => "00000000", 108 => "00010001", 109 => "11110111", 110 => "00010111", 111 => "00010100", 112 => "00001010", 113 => "00101001", 114 => "00011001", 115 => "00011101", 116 => "00101001", 117 => "00010110", 118 => "00000010", 119 => "00000001", 120 => "00000000", 121 => "01001101", 122 => "01000000", 123 => "00011000", 124 => "00000010", 125 => "00000000", 126 => "00001111", 127 => "00010011", 128 => "00011101", 129 => "00010011", 130 => "00101101", 131 => "00000010", 132 => "00000001", 133 => "00010010", 134 => "00001100", 135 => "01001101", 136 => "01000000", 137 => "00011000", 138 => "00000010", 139 => "00000011", 140 => "00000000", 141 => "00000011", 142 => "00010000", 143 => "00011010", 144 => "11011110", 145 => "00000010", 146 => "00000100", 147 => "00000111", 148 => "00000100", 149 => "00001011", 150 => "00001001", 151 => "00000011", 152 => "00001011", 153 => "01111001", 154 => "00000010", 155 => "00000110", 156 => "00000001", 157 => "00000111", 158 => "00000010", 159 => "00000001", 160 => "00000000", 161 => "00000011", 162 => "00010000", 163 => "00011010", 164 => "00010110", 165 => "00000101", 166 => "00011110", 167 => "00000000", 168 => "00010001", 169 => "11110111", 170 => "00010111", 171 => "00010100", 172 => "00001010", 173 => "00101001", 174 => "00011001", 175 => "00011101", 176 => "00101001", 177 => "00010110", 178 => "00000010", 179 => "00000001", 180 => "00000010", 181 => "01001101", 182 => "01000000", 183 => "00011000", 184 => "00000010", 185 => "00000000", 186 => "00001111", 187 => "00010011", 188 => "00011101", 189 => "00010011", 190 => "00101101", 191 => "00000010", 192 => "00010100", 193 => "00010010", 194 => "00001100", 195 => "00001100", 196 => "01000000", 197 => "00011000", 198 => "00000010", 199 => "00001100", 200 => "00000000", 201 => "00000011", 202 => "00010000", 203 => "00011010", 204 => "00010110", 205 => "00000000", 206 => "00001111", 207 => "00010011", 208 => "00011101", 209 => "00010011", 210 => "00101101", 211 => "00000010", 212 => "00010110", 213 => "00100010", 214 => "00001100", 215 => "00101011", 216 => "01000000", 217 => "00011000", 218 => "00000010", 219 => "00000001", 220 => "00000000", 221 => "00000011", 222 => "00010000", 223 => "00011010", 224 => "00010110", 225 => "00000000", 226 => "00001111", 227 => "00010011", 228 => "00011101", 229 => "00010011", 230 => "00101101", 231 => "00000010", 232 => "00010100", 233 => "00010010", 234 => "00001100", 235 => "01001101", 236 => "01000000", 237 => "00011000", 238 => "00000010", 239 => "00000001", 240 => "00000110", 241 => "00010011", 242 => "00101101", 243 => "00000010", 244 => "00010100", 245 => "00000001", 246 => "00001111", 247 => "00010011", 248 => "00011101", 249 => "00010011", 250 => "00101101", 251 => "00000010", 252 => "00010100", 253 => "00010010", 254 => "00001100", 255 => "00001100", 256 => "01000000", 257 => "00011000", 258 => "00000010", 259 => "00001100", 260 => "00000000", 261 => "00000011", 262 => "00010000", 263 => "00011010", 264 => "00010110", 265 => "11110101", 266 => "00001111", 267 => "00001101", 268 => "00000001", 269 => "00000001", 270 => "00000101", 271 => "00000011", 272 => "00000001", 273 => "00000001", 274 => "00000011", 275 => "00000101", 276 => "00000001", 277 => "00001001", 278 => "00000010", 279 => "00000001", 280 => "00000100", 281 => "00000011", 282 => "00000110", 283 => "00000110", 284 => "00010110", others => (others =>'0'));
                count <= 28;
            elsif count = 28 then
               --test # 28
                RAM <= (2 => "00010100", 3 => "00001110", 4 => "00010111",  5 => "00000001", 6 => "00010110", 7 => "00000001", 8 => "00000000", 9 => "00010100", 10 => "00000010", 11 => "00000010", 12 => "00000000", 13 => "00000011", 14 => "00001100", 15 => "00000010", 16 => "00000010", 17 => "00000001", 18 => "00010110", 19 => "00000001", 20 => "00000110", 21 => "01001101", 22 => "01000000", 23 => "00000010", 24 => "00000010", 25 => "00010101", 26 => "00000100", 27 => "00000111", 28 => "00000100", 29 => "00001011", 30 => "00001001", 31 => "00000011", 32 => "00001011", 33 => "01111001", 34 => "00000010", 35 => "00000110", 36 => "00000001", 37 => "00000111", 38 => "00000010", 39 => "00000001", 40 => "00000000", 41 => "00000011", 42 => "00010000", 43 => "00011010", 44 => "00010110", 45 => "00000110", 46 => "00000101", 47 => "10000010", 48 => "00001001", 49 => "10000100", 50 => "00001101", 51 => "00000011", 52 => "00010000", 53 => "00011010", 54 => "00010110", 55 => "00011010", 56 => "00011011", 57 => "00100010", 58 => "00000010", 59 => "00000011", 60 => "00000011", 61 => "01001101", 62 => "01000000", 63 => "00011000", 64 => "00000010", 65 => "00000110", 66 => "00001100", 67 => "00010010", 68 => "00000111", 69 => "10111110", 70 => "00000010", 71 => "00001111", 72 => "00001100", 73 => "00100111", 74 => "00010110", 75 => "00011100", 76 => "00001010", 77 => "00000000", 78 => "00000010", 79 => "00000001", 80 => "00000000", 81 => "00010011", 82 => "00101101", 83 => "00000010", 84 => "00010100", 85 => "00000101", 86 => "00011110", 87 => "00000000", 88 => "00010001", 89 => "11110111", 90 => "00010111", 91 => "00010100", 92 => "00001010", 93 => "00101001", 94 => "01000010", 95 => "00011101", 96 => "00101001", 97 => "00010110", 98 => "00000010", 99 => "00000001", 100 => "00000001", 101 => "00000011", 102 => "00010000", 103 => "00011010", 104 => "00010110", 105 => "00000101", 106 => "00011110", 107 => "00000000", 108 => "00010001", 109 => "11110111", 110 => "00010111", 111 => "00010100", 112 => "00001010", 113 => "00101001", 114 => "00011001", 115 => "00011101", 116 => "00101001", 117 => "00010110", 118 => "00000010", 119 => "00000001", 120 => "00000000", 121 => "01001101", 122 => "01000000", 123 => "00011000", 124 => "00000010", 125 => "00000000", 126 => "00001111", 127 => "00010011", 128 => "00011101", 129 => "00010011", 130 => "00101101", 131 => "00000010", 132 => "00000001", 133 => "00010010", 134 => "00001100", 135 => "01001101", 136 => "01000000", 137 => "00011000", 138 => "00000010", 139 => "00000011", 140 => "00000000", 141 => "00000011", 142 => "00010000", 143 => "00011010", 144 => "11011110", 145 => "00000010", 146 => "00000100", 147 => "00000111", 148 => "00000100", 149 => "00001011", 150 => "00001001", 151 => "00000011", 152 => "00001011", 153 => "01111001", 154 => "00000010", 155 => "00000110", 156 => "00000001", 157 => "00000111", 158 => "00000010", 159 => "00000001", 160 => "00000000", 161 => "00000011", 162 => "00010000", 163 => "00011010", 164 => "00010110", 165 => "00000101", 166 => "00011110", 167 => "00000000", 168 => "00010001", 169 => "11110111", 170 => "00010111", 171 => "00010100", 172 => "00001010", 173 => "00101001", 174 => "00011001", 175 => "00011101", 176 => "00101001", 177 => "00010110", 178 => "00000010", 179 => "00000001", 180 => "00000010", 181 => "01001101", 182 => "01000000", 183 => "00011000", 184 => "00000010", 185 => "00000000", 186 => "00001111", 187 => "00010011", 188 => "00011101", 189 => "00010011", 190 => "00101101", 191 => "00000010", 192 => "00010100", 193 => "00010010", 194 => "00001100", 195 => "00001100", 196 => "01000000", 197 => "00011000", 198 => "00000010", 199 => "00001100", 200 => "00000000", 201 => "00000011", 202 => "00010000", 203 => "00011010", 204 => "00010110", 205 => "00000000", 206 => "00001111", 207 => "00010011", 208 => "00011101", 209 => "00010011", 210 => "00101101", 211 => "00000010", 212 => "00010110", 213 => "00100010", 214 => "00001100", 215 => "00101011", 216 => "01000000", 217 => "00011000", 218 => "00000010", 219 => "00000001", 220 => "00000000", 221 => "00000011", 222 => "00010000", 223 => "00011010", 224 => "00010110", 225 => "00000000", 226 => "00001111", 227 => "00010011", 228 => "00011101", 229 => "00010011", 230 => "00101101", 231 => "00000010", 232 => "00010100", 233 => "00010010", 234 => "00001100", 235 => "01001101", 236 => "01000000", 237 => "00011000", 238 => "00000010", 239 => "00000001", 240 => "00000110", 241 => "00010011", 242 => "00101101", 243 => "00000010", 244 => "00010100", 245 => "00000001", 246 => "00001111", 247 => "00010011", 248 => "00011101", 249 => "00010011", 250 => "00101101", 251 => "00000010", 252 => "00010100", 253 => "00010010", 254 => "00001100", 255 => "00001100", 256 => "01000000", 257 => "00011000", 258 => "00000010", 259 => "00001100", 260 => "00000000", 261 => "00000011", 262 => "00010000", 263 => "00011010", 264 => "00010110", 265 => "00000010", 266 => "00001111", 267 => "00001101", 268 => "00000001", 269 => "00000001", 270 => "00000101", 271 => "00000011", 272 => "00000001", 273 => "00000001", 274 => "00000011", 275 => "00000101", 276 => "00000001", 277 => "00001001", 278 => "00000010", 279 => "00000001", 280 => "00000100", 281 => "00000011", 282 => "00000110", 283 => "00000110", 284 => "00010110", others => (others =>'0'));
                count <= 29;    
            elsif count = 29 then
               --test # 29
                RAM <= (2 => "00010100", 3 => "00001110", 4 => "01100101",  5 => "00000001", 6 => "00010110", 7 => "00000001", 8 => "00000000", 9 => "00010100", 10 => "00000010", 11 => "00000010", 12 => "00000000", 13 => "00000011", 14 => "00001100", 15 => "00000010", 16 => "00000010", 17 => "00000001", 18 => "00010110", 19 => "00000001", 20 => "00000110", 21 => "01001101", 22 => "01000000", 23 => "00000010", 24 => "00000010", 25 => "00010101", 26 => "00000100", 27 => "00000111", 28 => "00000100", 29 => "00001011", 30 => "00001001", 31 => "00000011", 32 => "00001011", 33 => "00001011", 34 => "00000010", 35 => "00000110", 36 => "00000001", 37 => "00000111", 38 => "00000010", 39 => "00000001", 40 => "00000000", 41 => "00000011", 42 => "00010000", 43 => "00011010", 44 => "00010110", 45 => "00000110", 46 => "00000101", 47 => "00001101", 48 => "00001001", 49 => "10000100", 50 => "00001101", 51 => "00000011", 52 => "00010000", 53 => "00011010", 54 => "00010110", 55 => "00011010", 56 => "00011011", 57 => "00100010", 58 => "00000010", 59 => "01110001", 60 => "00000011", 61 => "01001101", 62 => "01000000", 63 => "00011000", 64 => "00000010", 65 => "00000110", 66 => "00001100", 67 => "00010010", 68 => "00000111", 69 => "10111110", 70 => "00000010", 71 => "00001111", 72 => "00001100", 73 => "00100111", 74 => "00010110", 75 => "00011100", 76 => "00001010", 77 => "00000000", 78 => "00000010", 79 => "00000001", 80 => "00000000", 81 => "00010011", 82 => "00101101", 83 => "00000010", 84 => "00010100", 85 => "00000101", 86 => "00011110", 87 => "00000000", 88 => "00010001", 89 => "10010011", 90 => "00010111", 91 => "00010100", 92 => "00001010", 93 => "00101001", 94 => "01000010", 95 => "00011101", 96 => "00101001", 97 => "00010110", 98 => "00000010", 99 => "00000001", 100 => "00000001", 101 => "00000011", 102 => "00010000", 103 => "00011010", 104 => "00010110", 105 => "00000101", 106 => "00011110", 107 => "00000000", 108 => "00010001", 109 => "01101111", 110 => "00010111", 111 => "00010100", 112 => "00001010", 113 => "00101001", 114 => "00011001", 115 => "00011101", 116 => "00101001", 117 => "00010110", 118 => "00000010", 119 => "00000001", 120 => "00000000", 121 => "01001101", 122 => "01000000", 123 => "00011000", 124 => "00000010", 125 => "00000000", 126 => "00001111", 127 => "00010011", 128 => "00011101", 129 => "00010011", 130 => "00101101", 131 => "00000010", 132 => "00000001", 133 => "00010010", 134 => "00001100", 135 => "01001101", 136 => "01000000", 137 => "00011000", 138 => "00000010", 139 => "00000011", 140 => "00000000", 141 => "00000011", 142 => "00010000", 143 => "00011010", 144 => "00000010", 145 => "00000010", 146 => "00000100", 147 => "00000111", 148 => "00000100", 149 => "00001011", 150 => "00001001", 151 => "00000011", 152 => "00001011", 153 => "01111001", 154 => "00000010", 155 => "00000110", 156 => "00000001", 157 => "00000111", 158 => "00000010", 159 => "00000001", 160 => "00000000", 161 => "00000011", 162 => "00010000", 163 => "00011010", 164 => "00010110", 165 => "00000101", 166 => "00011110", 167 => "00000000", 168 => "00010001", 169 => "10010011", 170 => "00010111", 171 => "00010100", 172 => "00001010", 173 => "00101001", 174 => "00011001", 175 => "00011101", 176 => "00101001", 177 => "00010110", 178 => "00000010", 179 => "00000001", 180 => "00000010", 181 => "01001101", 182 => "01000000", 183 => "00011000", 184 => "00000010", 185 => "00000000", 186 => "00001111", 187 => "00010011", 188 => "00011101", 189 => "00010011", 190 => "00101101", 191 => "00000010", 192 => "00010100", 193 => "00010010", 194 => "00001100", 195 => "00001100", 196 => "01000000", 197 => "00011000", 198 => "00000010", 199 => "00001100", 200 => "00000000", 201 => "00000011", 202 => "00010000", 203 => "00011010", 204 => "00010110", 205 => "00000000", 206 => "00001111", 207 => "00010011", 208 => "00011101", 209 => "00010011", 210 => "00101101", 211 => "00000010", 212 => "00010110", 213 => "00100010", 214 => "00001100", 215 => "00101011", 216 => "01000000", 217 => "00011000", 218 => "00000010", 219 => "00000001", 220 => "00000000", 221 => "00000011", 222 => "00010000", 223 => "00011010", 224 => "00010110", 225 => "00000000", 226 => "00001111", 227 => "10111110", 228 => "00011101", 229 => "00010011", 230 => "00101101", 231 => "00000010", 232 => "00010100", 233 => "00010010", 234 => "00001100", 235 => "01001101", 236 => "10100100", 237 => "00011000", 238 => "00000010", 239 => "00000001", 240 => "00000110", 241 => "00010011", 242 => "00101101", 243 => "00000010", 244 => "00010100", 245 => "00000001", 246 => "00001111", 247 => "00010011", 248 => "00011101", 249 => "00010011", 250 => "00101101", 251 => "00000010", 252 => "00010100", 253 => "00010010", 254 => "00001100", 255 => "00001100", 256 => "01000000", 257 => "00011000", 258 => "00000010", 259 => "00001100", 260 => "00000000", 261 => "00000011", 262 => "00010000", 263 => "00011010", 264 => "00010110", 265 => "00000010", 266 => "00001111", 267 => "00001101", 268 => "00000001", 269 => "00000001", 270 => "00000101", 271 => "00000011", 272 => "00000001", 273 => "00000001", 274 => "00000011", 275 => "00000101", 276 => "00000001", 277 => "00001001", 278 => "00000010", 279 => "00000001", 280 => "00000100", 281 => "00000011", 282 => "00000110", 283 => "00000110", 284 => "00010110", others => (others =>'0'));
                count <= 30;
            elsif count = 30 then
               --test # 30
                RAM <= (2 => "00010100", 3 => "00001110", 4 => "00011111",  5 => "00000001", 6 => "00010110", 7 => "00000001", 8 => "00000000", 9 => "00010100", 10 => "00000010", 11 => "00000010", 12 => "00000000", 13 => "00000011", 14 => "00001100", 15 => "00000010", 16 => "00000010", 17 => "00000001", 18 => "00010110", 19 => "00000001", 20 => "00000110", 21 => "01001101", 22 => "01000000", 23 => "00000010", 24 => "00000010", 25 => "00010101", 26 => "00000100", 27 => "00000111", 28 => "00000100", 29 => "00001011", 30 => "00001001", 31 => "00000011", 32 => "00001011", 33 => "00001011", 34 => "00000010", 35 => "00000110", 36 => "00000001", 37 => "00000111", 38 => "00000010", 39 => "00000001", 40 => "00000000", 41 => "00000011", 42 => "00010000", 43 => "00011010", 44 => "00010110", 45 => "00000110", 46 => "00000101", 47 => "00001101", 48 => "00001001", 49 => "10000100", 50 => "00001101", 51 => "00000011", 52 => "00010000", 53 => "00011010", 54 => "00010110", 55 => "00011010", 56 => "00011011", 57 => "00100010", 58 => "00000010", 59 => "01110001", 60 => "00000011", 61 => "01001101", 62 => "01000000", 63 => "00011000", 64 => "00000010", 65 => "00000110", 66 => "00001100", 67 => "00010010", 68 => "00000111", 69 => "10111110", 70 => "00000010", 71 => "00001111", 72 => "00001100", 73 => "00100111", 74 => "00010110", 75 => "00011100", 76 => "00001010", 77 => "00000000", 78 => "00000010", 79 => "00000001", 80 => "00000000", 81 => "00010011", 82 => "00101101", 83 => "00000010", 84 => "00010100", 85 => "00000101", 86 => "00011110", 87 => "00000000", 88 => "00010001", 89 => "10010011", 90 => "00010111", 91 => "00010100", 92 => "00001010", 93 => "00101001", 94 => "01000010", 95 => "00011101", 96 => "00101001", 97 => "00010110", 98 => "00000010", 99 => "00000001", 100 => "00000001", 101 => "00000011", 102 => "00010000", 103 => "00011010", 104 => "00010110", 105 => "00000101", 106 => "00011110", 107 => "00000000", 108 => "00010001", 109 => "01101111", 110 => "00010111", 111 => "00010100", 112 => "00001010", 113 => "00101001", 114 => "00011001", 115 => "00011101", 116 => "00101001", 117 => "00010110", 118 => "00000010", 119 => "00000001", 120 => "00000000", 121 => "01001101", 122 => "01000000", 123 => "00011000", 124 => "00000010", 125 => "00000000", 126 => "00001111", 127 => "00010011", 128 => "00011101", 129 => "00010011", 130 => "00101101", 131 => "00000010", 132 => "00000001", 133 => "00010010", 134 => "00001100", 135 => "01001101", 136 => "01000000", 137 => "00011000", 138 => "00000010", 139 => "00000011", 140 => "00000000", 141 => "00000011", 142 => "00010000", 143 => "00011010", 144 => "00000010", 145 => "00000010", 146 => "00000100", 147 => "00000111", 148 => "00000100", 149 => "00001011", 150 => "00001001", 151 => "00000011", 152 => "00001011", 153 => "01111001", 154 => "00000010", 155 => "00000110", 156 => "00000001", 157 => "00000111", 158 => "00000010", 159 => "00000001", 160 => "00000000", 161 => "00000011", 162 => "00010000", 163 => "00011010", 164 => "00010110", 165 => "00000101", 166 => "00011110", 167 => "00000000", 168 => "00010001", 169 => "10010011", 170 => "00010111", 171 => "00010100", 172 => "00001010", 173 => "00101001", 174 => "00011001", 175 => "00011101", 176 => "00101001", 177 => "00010110", 178 => "00000010", 179 => "00000001", 180 => "00000010", 181 => "01001101", 182 => "01000000", 183 => "00011000", 184 => "00000010", 185 => "00000000", 186 => "00001111", 187 => "00010011", 188 => "00011101", 189 => "00010011", 190 => "00101101", 191 => "00000010", 192 => "00010100", 193 => "00010010", 194 => "00001100", 195 => "00001100", 196 => "01000000", 197 => "00011000", 198 => "00000010", 199 => "00001100", 200 => "00000000", 201 => "00000011", 202 => "00010000", 203 => "00011010", 204 => "00010110", 205 => "00000000", 206 => "00001111", 207 => "00010011", 208 => "00011101", 209 => "00010011", 210 => "00101101", 211 => "00000010", 212 => "00010110", 213 => "00100010", 214 => "00001100", 215 => "00101011", 216 => "01000000", 217 => "00011000", 218 => "00000010", 219 => "00000001", 220 => "00000000", 221 => "00000011", 222 => "00010000", 223 => "00011010", 224 => "00010110", 225 => "00000000", 226 => "00001111", 227 => "10111110", 228 => "00011101", 229 => "00010011", 230 => "00101101", 231 => "00000010", 232 => "00010100", 233 => "00010010", 234 => "00001100", 235 => "01001101", 236 => "10100100", 237 => "00011000", 238 => "00000010", 239 => "00000001", 240 => "00000110", 241 => "00010011", 242 => "00101101", 243 => "00000010", 244 => "00010100", 245 => "00000001", 246 => "00001111", 247 => "00010011", 248 => "00011101", 249 => "00010011", 250 => "00101101", 251 => "00000010", 252 => "00010100", 253 => "00010010", 254 => "00001100", 255 => "00001100", 256 => "01000000", 257 => "00011000", 258 => "00000010", 259 => "00001100", 260 => "00000000", 261 => "00000011", 262 => "00010000", 263 => "00011010", 264 => "00010110", 265 => "00000010", 266 => "00001111", 267 => "00001101", 268 => "00000001", 269 => "00000001", 270 => "00000101", 271 => "00000011", 272 => "00000001", 273 => "00000001", 274 => "00000011", 275 => "00000101", 276 => "00000001", 277 => "00001001", 278 => "00000010", 279 => "00000001", 280 => "00000100", 281 => "00000011", 282 => "00000110", 283 => "00000110", 284 => "00010110", others => (others =>'0'));
                count<=31;
            elsif count=31 then
                --test #31
                RAM <= (2 => "11111111", 3 =>"11111111",4 => "00000001", 30 => "00000011", 31 => "00000011", 32 => "00000011", 33 => "00000011", 36 => "00000111", 259=>"11111111", 285 =>"00001000" , 291 =>"00001000" ,600=>"11111111",others => (others =>'0'));
                count<=32;
            elsif count=32 then
                --test #32
                
               RAM <= (2 => "11111111", 3 =>"11111111",4 => "00000001", 5=>"11111111", 30 => "00000011", 31 => "00000011", 32 => "00000011", 33 => "00000011", 36 => "00000111", 259=>"11111111", 285 =>"00001000" , 291 =>"00001000" ,600=>"11111111",65029=>"11111111",65030=>"11101111", 65031=>"11110011",others => (others =>'1'));
               count<=33;
            elsif count=33 then
               --test #33
               RAM <= (2 => "00000100", 3 =>"00000101",4 => "00000011", 5=>"11111111", 20=>"00001111", 24=>"01010111", 25=>"00111111",26=>"00011111", 27=>"11111111", 30 => "00000011", 31 => "00000011", 32 => "00000011", 33 => "00000011", 36 => "00000111", 259=>"11111111", 285 =>"00001000" , 291 =>"00001000" ,600=>"11111111",65029=>"11111111",65030=>"11101111", 65031=>"11110011",others => (others =>'0'));
               count<=34;
            elsif count=34 then
               --test #34
               RAM <= (2 => "11111111", 3 =>"11111111",4 => "00000001", 654=>"01111111",others => (others =>'0'));
               count<=35;
            elsif count=35 then
               --test #35
               RAM <= (2 => "11111111", 3 =>"11111111",4 => "00000001", 5=>"01111111",others => (others =>'0'));
               count<=36;
            elsif count=36 then
                --test #36
                RAM <= (2 => "11111111", 3 =>"11111111",4 => "00000001", 65029=>"01111111",others => (others =>'0'));
                count<=37;
            elsif count=37 then
                --test #37
                RAM <= (2 => "00000100", 3 =>"00000101",4 => "00000011", 6=>"11111111", 7=>"00001111", 9=>"01010111", 15=>"00111111",23=>"00011111", 27=>"11111111", 30 => "00000011", 31 => "00000011", 32 => "00000011", 33 => "00000011", 36 => "00000111", 259=>"11111111", 285 =>"00001000" , 291 =>"00001000" ,600=>"11111111",65029=>"11111111",65030=>"11101111", 65031=>"11110011",others => (others =>'0'));
                count<=38;
            elsif count<=38 then
                --test #38
                RAM <= (2 => "00001000", 3 =>"00000111",4 => "00000011", 19=>"11111111", 24=>"00001111", 46=>"01010111", 60=>"00111111",others => (others =>'0'));
                count<=39;
            elsif count<=39 then
               --test #39
               RAM <= (2 => "00001000", 3 =>"00000111",4 => "00000011", 5=>"11001100", 12=>"11000111",19=>"11111111", 24=>"00001111", 46=>"01010111", 60=>"00111111",others => (others =>'0'));
                count<=40;
            elsif count=40 then
                --test #40
               RAM <= (2 => "00010100", 3 =>"00010000",4 => "00000011", 6=>"11001100", 13=>"11000111",17=>"11111111", 31=>"00001111", 97=>"01010111", 103=>"00111111",118=>"11111111", 131=>"00001111", 190=>"01010111", 217=>"00111111",284=>"00111111", others => (others =>'0'));
                count<=41;
            elsif count=41 then
               --test #41
               RAM <= (2 => "00001000", 3 =>"00000111",4 => "00000011", 16=>"11001100", 32=>"11000111",others => (others =>'0'));
               count<=42;
            elsif count=42 then
              --test #42
              RAM <= (2 => "00001000", 3 =>"00000111",4 => "00000011", 16=>"11001100", 19=>"11000111",others => (others =>'0'));
              count<=43;
            elsif count=43 then
              --test #43
              RAM <= (2 => "00000000", 3 => "00000000", 4 => "11111010",  5 => "00001101", 6 => "00000010", 7 => "00000001", 8 => "00000000", 9 => "00010100", 10 => "00000010", 11 => "00000010", 12 => "00000000", 13 => "00000011", 14 => "00001100", 15 => "00000010", 16 => "00000010", 17 => "00000001", 18 => "00010110", 19 => "00000001", 20 => "00000000", 21 => "00000010", 22 => "00000100", 23 => "00000111", 24 => "00000100", 25 => "00001011", 26 => "00001001", 27 => "00000011", 28 => "00001011", 29 => "01111001", 30 => "00000010", 31 => "00000110", 32 => "00000001", 33 => "00000111", 34 => "00000010", 35 => "00000001", 36 => "00000000", 37 => "00000110", 38 => "00000101", 39 => "10000010", 40 => "00001001", 41 => "10000100", 42 => "00001101", 43 => "00000011", 44 => "00010000", 45 => "00011010", 46 => "00010110", 47 => "00011010", 48 => "00011011", 49 => "00100010", 50 => "00000010", 51 => "00000011", 52 => "00000000", 53 => "00000110", 54 => "00001100", 55 => "00010010", 56 => "00000111", 57 => "10111110", 58 => "00000010", 59 => "00001111", 60 => "00001100", 61 => "00100111", 62 => "00010110", 63 => "00011100", 64 => "00001010", 65 => "00000000", 66 => "00000010", 67 => "00000001", 68 => "00000000", 69 => "00000101", 70 => "00011110", 71 => "00000000", 72 => "00010001", 73 => "11110111", 74 => "00010111", 75 => "00010100", 76 => "00001010", 77 => "00101001", 78 => "00011001", 79 => "00011101", 80 => "00101001", 81 => "00010110", 82 => "00000010", 83 => "00000001", 84 => "00000000", 85 => "00001010", 86 => "00001100", 87 => "00001101", 88 => "00010101", 89 => "00010110", 90 => "11100111", 91 => "10011011", 92 => "00000000", 93 => "00001010", 94 => "00010001", 95 => "00011001", 96 => "00001101", 97 => "00110010", 98 => "00000010", 99 => "00000001", 100 => "00000100", 101 => "00000000", 102 => "00001111", 103 => "00010011", 104 => "00011101", 105 => "00010011", 106 => "00101101", 107 => "00000010", 108 => "00010100", 109 => "00010010", 110 => "00001100", 111 => "01001101", 112 => "01000000", 113 => "00011000", 114 => "00000010", 115 => "00000011", 116 => "00000000", 117 => "00000000", 118 => "00001111", 119 => "00010011", 120 => "00011101", 121 => "00010011", 122 => "00101101", 123 => "00000010", 124 => "00010100", 125 => "00100010", 126 => "00001100", 127 => "01001101", 128 => "01000000", 129 => "00011000", 130 => "00000010", 131 => "00000001", 132 => "00000000", 133 => "00000000", 134 => "00001111", 135 => "00010011", 136 => "00011101", 137 => "00010011", 138 => "00101101", 139 => "00000010", 140 => "00010100", 141 => "00010010", 142 => "00001100", 143 => "01001101", 144 => "01000000", 145 => "00011000", 146 => "00000010", 147 => "00000001", 148 => "00000110", 149 => "00000000", 150 => "00001111", 151 => "00010011", 152 => "00011101", 153 => "00010011", 154 => "00101101", 155 => "00000010", 156 => "00010100", 157 => "00010010", 158 => "00001100", 159 => "01001101", 160 => "01000000", 161 => "00011000", 162 => "00000010", 163 => "00001100", 164 => "00000000", 165 => "00001101", 166 => "00010000", 167 => "00001101", 168 => "10000110", 169 => "00000001", 170 => "00000101", 171 => "00111111", 172 => "00000001", 173 => "00011111", 174 => "00111111", 175 => "00101101", 176 => "00010101", 177 => "00001001", 178 => "00000010", 179 => "00000001", 180 => "00000000", others => (others =>'0'));
              count<=44;
            elsif count=44 then
              --test #44
              RAM <= (2 => "11110111", 3 =>"11011111",4 => "00000101", 654=>"01111111",others => (others =>'0'));
              count<=45;
            elsif count=45 then
              --test #45
              RAM <= (2 => "00000001", 3 =>"00000001",4 => "00000101", 5=>"01111111",others => (others =>'0'));
              count<=46;
            elsif count=46 then
              --test #46
              RAM <= (2 => "11111111", 3 =>"11111111",4 => "00000001", 65000=>"01111111",others => (others =>'0'));
              count<=47;
            elsif count=47 then
              --test #47
              RAM <= (2 => "11111111", 3 =>"11111111",4 => "00000001", 260=>"01111111",others => (others =>'0'));
              count<=48;
            elsif count=48 then
              --test #48
              RAM <= (2 => "00001000", 3 =>"00000111",4 => "00000011", 12=>"11001100", 28=>"11000111",52=>"11111111", others => (others =>'0'));
              count<=49;
            elsif count=49 then
               --test #49 FEDE prima riga completa
               RAM <= (2 => "10000000", 3 =>"10000000",4 => "01000000", 5=>"11001100", 132=>"11000111", others => (others =>'0'));
               count<=50;
            elsif count=50 then
                --test #50 FEDE ultima riga completa
                RAM <= (2 => "10000000", 3 =>"10000000",4 => "01000000", 16261=>"11001100", 16388=>"11000111", others => (others =>'0'));
                count<=51;             
             elsif count=51 then
                --test #51 FEDE prima colonna completa
                RAM <= (2 => "10000000", 3 =>"10000000",4 => "01000000", 5=>"11001100", 16261=>"11000111", others => (others =>'0'));
                count<=52;
             elsif count=52 then
                --test #52 FEDE ultima colonna completa
               RAM <= (2 => "10000000", 3 =>"10000000",4 => "01000000", 132=>"11001100", 16388=>"11000111", others => (others =>'0'));
               count<=53;
            elsif count=53 then
                --test #53 FEDE quadratino 2x2 in centro
                RAM <= (2 => "10000000", 3 =>"10000000",4 => "01000000", 12168=>"11001100", 12169=>"11001100",12296=>"11001100", 12297=>"11001100", others => (others =>'0'));
                count<=54;
            
            elsif count=54 then
                --test #54 FEDE tutta piena
                RAM <= (2 => "11111111", 3 =>"11111111",4 => "01000000", others => ("11111111"));
                count<=55;
                
            elsif count = 55 then
                --test #55 SERGIO E MARCO prima casella inferiore alla soglia, tutto il resto maggiore della soglia
                RAM <= (2 => "11111111", 3 =>"11111111", 4 => "10000000", 5 => "01111111", others => ("10000001"));     
                count<=56;
                
            elsif count = 56 then
                --test #56 SERGIO E MARCO prima casella inferiore alla soglia, tutto il resto uguale alla soglia
                RAM <= (2 => "11111111", 3 =>"11111111", 4 => "10000000", 5 => "01111111", others => ("10000000"));
                count<=57;
                
            elsif count = 57 then
                --test #57 SERGIO E MARCO matrice 4x4 con 1� riga e 1� colonna superiori alla soglia, il resto inferiore
                RAM <= (2 => "00000100", 3 => "00000100", 4 => "00000001", 5 => "00000010", 6 => "00000010", 7 => "00000010", 8 => "00000010", 9 => "00000010", 13 => "00000010", 17 => "00000010", others => (others =>'0'));        
                count<=58;
                
            elsif count = 58 then
                --test #58 SERGIO E MARCO matrice 4x4 con 1� riga e 1� colonna inferiori alla soglia, il resto superiore
                RAM <= (2 => "00000100", 3 => "00000100", 4 => "00000011", 5 => "00000010", 6 => "00000010", 7 => "00000010", 8 => "00000010", 9 => "00000010", 13 => "00000010", 17 => "00000010", others => ("00000101"));        
                count<=59;
                
           elsif count = 59 then
               --test #59 SERGIO E MARCO matrice 4x4 con due soli valori sopra la soglia (1x2 e 3x3)
               RAM <= (2 => "00000100", 3 => "00000100", 4 => "00000001", 6 => "00000010", 13 => "00000010", others => (others =>'0'));
               count<=60;
               
          elsif count = 60 then
              --test #60 SERGIO E MARCO matrice 4x4 con il solo valore in basso a dx maggiore della soglia
              RAM <= (2 => "00000100", 3 => "00000100", 4 => "00000001", 20 => "00000010", others => (others =>'0'));
              count<=61;  
         
          elsif count = 61 then
              --test #61 SERGIO E MARCO matrice 4x4 con il solo valore in basso a dx minore della soglia
              RAM <= (2 => "00000100", 3 => "00000100", 4 => "00000001", 20 => "00000000", others => ("11111111"));
              count<=62;
              
          elsif count = 62 then
              --test #62 SERGIO E MARCO matrice 1x1 con valore minore della soglia
              RAM <= (2 => "00000001", 3 => "00000001", 4 => "00000001", 5 => "00000000", others => ("00000000"));
              count<=63;  
              
          elsif count = 63 then
                  --test #63 SERGIO E MARCO matrice 1x1 con valore maggiore della soglia
                  RAM <= (2 => "00000001", 3 => "00000001", 4 => "00000001", 5 => "00000100", others => ("00000000"));
                  count<=64;
                    
          elsif count = 64 then
                  --test #64 SERGIO E MARCO matrice 4x4 con tre valori maggiori della soglia (2x1, 2x4, 4x2)
                  RAM <= (2 => "00000100", 3 => "00000100", 4 => "00000001", 9 => "00000100", 12 => "00000100", 18 => "00000100", others => (others =>'0'));
                  count<=65;
                  
          elsif count = 65 then
                  --test #65 SERGIO E MARCO matrice 4x4 con due valori maggiori della soglia (4x1, 3x2)
                  RAM <= (2 => "00000100", 3 => "00000100", 4 => "00000001", 14 => "00000100", 17 => "00000100", others => (others =>'0'));
                  count<=66;                                                              
                       
            end if;   
               
          else
             mem_o_data <= RAM(conv_integer(mem_address)) after 1 ns;   
          end if;
      end if;
     end if;
    end if;
   end process;
 
  
test : process is
begin 

        --test # 0
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);

        assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
        assert RAM(0) = "00010101" report "FAIL low bits" severity failure;

        --test # 1
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);

        assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
        assert RAM(0) = "10101000" report "FAIL low bits" severity failure;


        --test # 2
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);

        assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
        assert RAM(0) = "00000000" report "FAIL low bits" severity failure;


        --test # 3
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);

        assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
        assert RAM(0) = "00000000" report "FAIL low bits" severity failure;

        
        --test # 4
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);

        assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
        assert RAM(0) = "00000000" report "FAIL low bits" severity failure;

        
        --test # 5
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);

        assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
        assert RAM(0) = "00000001" report "FAIL low bits" severity failure;
        
        
        --test # 6
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);

        assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
        assert RAM(0) = "00000001" report "FAIL low bits" severity failure;
        
        --test # 7
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);

        assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
        assert RAM(0) = "00000001" report "FAIL low bits" severity failure;
        
        --test # 8
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);

        assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
        assert RAM(0) = "00000110" report "FAIL low bits" severity failure;
        
        
        --test # 9
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);

        assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
        assert RAM(0) = "00000100" report "FAIL low bits" severity failure;
        
        --test # 10
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);

        assert RAM(1) = "11111110" report "FAIL high bits" severity failure;
        assert RAM(0) = "00000001" report "FAIL low bits" severity failure;
        
        
        --test # 11
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);

        assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
        assert RAM(0) = "00000000" report "FAIL low bits" severity failure;
     
        
        --test # 12
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);

        assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
        assert RAM(0) = "00110110" report "FAIL low bits" severity failure;
        
        --test # 13
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);

        assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
        assert RAM(0) = "00000001" report "FAIL low bits" severity failure;
        
        --test # 14
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);

        assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
        assert RAM(0) = "00001110" report "FAIL low bits" severity failure;
        
        --test # 15
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);

        assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
        assert RAM(0) = "00001000" report "FAIL low bits" severity failure;
        
        --test # 16
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);

        assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
        assert RAM(0) = "00011110" report "FAIL low bits" severity failure;
        
        --test # 17
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);

        assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
        assert RAM(0) = "01001101" report "FAIL low bits" severity failure;
        
        --test # 18
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);

        assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
        assert RAM(0) = "00101010" report "FAIL low bits" severity failure;
        
        --test # 19
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);

        assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
        assert RAM(0) = "01010100" report "FAIL low bits" severity failure;
        
        --test # 20
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);

        assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
        assert RAM(0) = "00000100" report "FAIL low bits" severity failure;
        
        --test # 21
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);

        assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
        assert RAM(0) = "10100101" report "FAIL low bits" severity failure;
        
        --test # 22
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);

        assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
        assert RAM(0) = "00101101" report "FAIL low bits" severity failure;
        
        --test # 23
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);

        assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
        assert RAM(0) = "00000000" report "FAIL low bits" severity failure;
        
        --test # 24
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);

        assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
        assert RAM(0) = "00010000" report "FAIL low bits" severity failure;
        
        --test # 25
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);

        assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
        assert RAM(0) = "00000010" report "FAIL low bits" severity failure;
        
        --test # 26
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);

        assert RAM(1) = "00000001" report "FAIL high bits" severity failure;
        assert RAM(0) = "00001010" report "FAIL low bits" severity failure;
        
        --test # 27
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);

        assert RAM(1) = "00000001" report "FAIL high bits" severity failure;
        assert RAM(0) = "00011000" report "FAIL low bits" severity failure;
        
        --test # 28
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);

        assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
        assert RAM(0) = "11110111" report "FAIL low bits" severity failure;
        
        --test # 29
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);

        assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
        assert RAM(0) = "10000010" report "FAIL low bits" severity failure;
        
        --test # 30
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);

        assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
        assert RAM(0) = "11010000" report "FAIL low bits" severity failure;
        
        --test # 31
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);

        assert RAM(1) = "00000010" report "FAIL high bits" severity failure;
        assert RAM(0) = "10110010" report "FAIL low bits" severity failure;
        
        --test # 32
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);

        assert RAM(1) = "11111110" report "FAIL high bits" severity failure;
        assert RAM(0) = "00000001" report "FAIL low bits" severity failure;
        
         --test # 33
       wait for 100 ns;
       wait for c_CLOCK_PERIOD;
       tb_rst <= '1';
       wait for c_CLOCK_PERIOD;
       tb_rst <= '0';
       wait for c_CLOCK_PERIOD;
       tb_start <= '1';
       wait for c_CLOCK_PERIOD;
       tb_start <= '0';
       wait until tb_done = '1';
       wait until tb_done = '0';
       wait until rising_edge(tb_clk);

       assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
       assert RAM(0) = "00010100" report "FAIL low bits" severity failure;
       
          --test # 34
       wait for 100 ns;
       wait for c_CLOCK_PERIOD;
       tb_rst <= '1';
       wait for c_CLOCK_PERIOD;
       tb_rst <= '0';
       wait for c_CLOCK_PERIOD;
       tb_start <= '1';
       wait for c_CLOCK_PERIOD;
       tb_start <= '0';
       wait until tb_done = '1';
       wait until tb_done = '0';
       wait until rising_edge(tb_clk);

       assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
       assert RAM(0) = "00000001" report "FAIL low bits" severity failure;
       --test # 35
       wait for 100 ns;
       wait for c_CLOCK_PERIOD;
       tb_rst <= '1';
       wait for c_CLOCK_PERIOD;
       tb_rst <= '0';
       wait for c_CLOCK_PERIOD;
       tb_start <= '1';
       wait for c_CLOCK_PERIOD;
       tb_start <= '0';
       wait until tb_done = '1';
       wait until tb_done = '0';
       wait until rising_edge(tb_clk);

       assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
       assert RAM(0) = "00000001" report "FAIL low bits" severity failure;
       --test # 36
       wait for 100 ns;
       wait for c_CLOCK_PERIOD;
       tb_rst <= '1';
       wait for c_CLOCK_PERIOD;
       tb_rst <= '0';
       wait for c_CLOCK_PERIOD;
       tb_start <= '1';
       wait for c_CLOCK_PERIOD;
       tb_start <= '0';
       wait until tb_done = '1';
       wait until tb_done = '0';
       wait until rising_edge(tb_clk);

       assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
       assert RAM(0) = "00000001" report "FAIL low bits" severity failure;
       
        --test # 37
         wait for 100 ns;
         wait for c_CLOCK_PERIOD;
         tb_rst <= '1';
         wait for c_CLOCK_PERIOD;
         tb_rst <= '0';
         wait for c_CLOCK_PERIOD;
         tb_start <= '1';
         wait for c_CLOCK_PERIOD;
         tb_start <= '0';
         wait until tb_done = '1';
         wait until tb_done = '0';
         wait until rising_edge(tb_clk);
    
         assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
         assert RAM(0) = "00001111" report "FAIL low bits" severity failure;
         
         
         --test # 38
          wait for 100 ns;
          wait for c_CLOCK_PERIOD;
          tb_rst <= '1';
          wait for c_CLOCK_PERIOD;
          tb_rst <= '0';
          wait for c_CLOCK_PERIOD;
          tb_start <= '1';
          wait for c_CLOCK_PERIOD;
          tb_start <= '0';
          wait until tb_done = '1';
          wait until tb_done = '0';
          wait until rising_edge(tb_clk);
     
          assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
          assert RAM(0) = "00101010" report "FAIL low bits" severity failure;
          
        --test # 39
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);
   
        assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
        assert RAM(0) = "00111000" report "FAIL low bits" severity failure;
        
        --test #40
        wait for 100 ns;
        wait for c_CLOCK_PERIOD;
        tb_rst <= '1';
        wait for c_CLOCK_PERIOD;
        tb_rst <= '0';
        wait for c_CLOCK_PERIOD;
        tb_start <= '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '1';
        wait until tb_done = '0';
        wait until rising_edge(tb_clk);
   
        assert RAM(1) = "00000001" report "FAIL high bits" severity failure;
        assert RAM(0) = "00001010" report "FAIL low bits" severity failure;
        
       --test #41
       wait for 100 ns;
       wait for c_CLOCK_PERIOD;
       tb_rst <= '1';
       wait for c_CLOCK_PERIOD;
       tb_rst <= '0';
       wait for c_CLOCK_PERIOD;
       tb_start <= '1';
       wait for c_CLOCK_PERIOD;
       tb_start <= '0';
       wait until tb_done = '1';
       wait until tb_done = '0';
       wait until rising_edge(tb_clk);
  
       assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
       assert RAM(0) = "00000011" report "FAIL low bits" severity failure;
       
       --test #42
      wait for 100 ns;
      wait for c_CLOCK_PERIOD;
      tb_rst <= '1';
      wait for c_CLOCK_PERIOD;
      tb_rst <= '0';
      wait for c_CLOCK_PERIOD;
      tb_start <= '1';
      wait for c_CLOCK_PERIOD;
      tb_start <= '0';
      wait until tb_done = '1';
      wait until tb_done = '0';
      wait until rising_edge(tb_clk);
 
      assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
      assert RAM(0) = "00000100" report "FAIL low bits" severity failure;
      
        --test #43
      wait for 100 ns;
      wait for c_CLOCK_PERIOD;
      tb_rst <= '1';
      wait for c_CLOCK_PERIOD;
      tb_rst <= '0';
      wait for c_CLOCK_PERIOD;
      tb_start <= '1';
      wait for c_CLOCK_PERIOD;
      tb_start <= '0';
      wait until tb_done = '1';
      wait until tb_done = '0';
      wait until rising_edge(tb_clk);
 
      assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
      assert RAM(0) = "00000000" report "FAIL low bits" severity failure;
      
      --test #44
      wait for 100 ns;
     wait for c_CLOCK_PERIOD;
     tb_rst <= '1';
     wait for c_CLOCK_PERIOD;
     tb_rst <= '0';
     wait for c_CLOCK_PERIOD;
     tb_start <= '1';
     wait for c_CLOCK_PERIOD;
     tb_start <= '0';
     wait until tb_done = '1';
     wait until tb_done = '0';
     wait until rising_edge(tb_clk);

     assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
     assert RAM(0) = "00000001" report "FAIL low bits" severity failure;
     
     --test #45
      wait for 100 ns;
     wait for c_CLOCK_PERIOD;
     tb_rst <= '1';
     wait for c_CLOCK_PERIOD;
     tb_rst <= '0';
     wait for c_CLOCK_PERIOD;
     tb_start <= '1';
     wait for c_CLOCK_PERIOD;
     tb_start <= '0';
     wait until tb_done = '1';
     wait until tb_done = '0';
     wait until rising_edge(tb_clk);

     assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
     assert RAM(0) = "00000001" report "FAIL low bits" severity failure;
     
       --test #46
       wait for 100 ns;
      wait for c_CLOCK_PERIOD;
      tb_rst <= '1';
      wait for c_CLOCK_PERIOD;
      tb_rst <= '0';
      wait for c_CLOCK_PERIOD;
      tb_start <= '1';
      wait for c_CLOCK_PERIOD;
      tb_start <= '0';
      wait until tb_done = '1';
      wait until tb_done = '0';
      wait until rising_edge(tb_clk);
 
      assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
      assert RAM(0) = "00000001" report "FAIL low bits" severity failure;
      
        --test #47
        wait for 100 ns;
       wait for c_CLOCK_PERIOD;
       tb_rst <= '1';
       wait for c_CLOCK_PERIOD;
       tb_rst <= '0';
       wait for c_CLOCK_PERIOD;
       tb_start <= '1';
       wait for c_CLOCK_PERIOD;
       tb_start <= '0';
       wait until tb_done = '1';
       wait until tb_done = '0';
       wait until rising_edge(tb_clk);
  
       assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
       assert RAM(0) = "00000001" report "FAIL low bits" severity failure;
       
      --test #48
      wait for 100 ns;
     wait for c_CLOCK_PERIOD;
     tb_rst <= '1';
     wait for c_CLOCK_PERIOD;
     tb_rst <= '0';
     wait for c_CLOCK_PERIOD;
     tb_start <= '1';
     wait for c_CLOCK_PERIOD;
     tb_start <= '0';
     wait until tb_done = '1';
     wait until tb_done = '0';
     wait until rising_edge(tb_clk);

     assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
     assert RAM(0) = "00000110" report "FAIL low bits" severity failure;

   --test #49
     wait for 100 ns;
     wait for c_CLOCK_PERIOD;
     tb_rst <= '1';
     wait for c_CLOCK_PERIOD;
     tb_rst <= '0';
     wait for c_CLOCK_PERIOD;
     tb_start <= '1';
     wait for c_CLOCK_PERIOD;
     tb_start <= '0';
     wait until tb_done = '1';
     wait until tb_done = '0';
     wait until rising_edge(tb_clk);

     assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
     assert RAM(0) = "10000000" report "FAIL low bits" severity failure;
     
      --test #50
          wait for 100 ns;
          wait for c_CLOCK_PERIOD;
          tb_rst <= '1';
          wait for c_CLOCK_PERIOD;
          tb_rst <= '0';
          wait for c_CLOCK_PERIOD;
          tb_start <= '1';
          wait for c_CLOCK_PERIOD;
          tb_start <= '0';
          wait until tb_done = '1';
          wait until tb_done = '0';
          wait until rising_edge(tb_clk);
     
          assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
          assert RAM(0) = "10000000" report "FAIL low bits" severity failure;
      --test #51
          wait for 100 ns;
          wait for c_CLOCK_PERIOD;
          tb_rst <= '1';
          wait for c_CLOCK_PERIOD;
          tb_rst <= '0';
          wait for c_CLOCK_PERIOD;
          tb_start <= '1';
          wait for c_CLOCK_PERIOD;
          tb_start <= '0';
          wait until tb_done = '1';
          wait until tb_done = '0';
          wait until rising_edge(tb_clk);
              
          assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
          assert RAM(0) = "10000000" report "FAIL low bits" severity failure;
    --test #52
          wait for 100 ns;
          wait for c_CLOCK_PERIOD;
          tb_rst <= '1';
          wait for c_CLOCK_PERIOD;
          tb_rst <= '0';
          wait for c_CLOCK_PERIOD;
          tb_start <= '1';
          wait for c_CLOCK_PERIOD;
          tb_start <= '0';
          wait until tb_done = '1';
          wait until tb_done = '0';
          wait until rising_edge(tb_clk);
                       
          assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
          assert RAM(0) = "10000000" report "FAIL low bits" severity failure;

    --test #53
          wait for 100 ns;
          wait for c_CLOCK_PERIOD;
          tb_rst <= '1';
          wait for c_CLOCK_PERIOD;
          tb_rst <= '0';
          wait for c_CLOCK_PERIOD;
          tb_start <= '1';
          wait for c_CLOCK_PERIOD;
          tb_start <= '0';
          wait until tb_done = '1';
          wait until tb_done = '0';
          wait until rising_edge(tb_clk);
                       
          assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
          assert RAM(0) = "00000100" report "FAIL low bits" severity failure;



    --test #54
          wait for 100 ns;
          wait for c_CLOCK_PERIOD;
          tb_rst <= '1';
          wait for c_CLOCK_PERIOD;
          tb_rst <= '0';
          wait for c_CLOCK_PERIOD;
          tb_start <= '1';
          wait for c_CLOCK_PERIOD;
          tb_start <= '0';
          wait until tb_done = '1';
          wait until tb_done = '0';
          wait until rising_edge(tb_clk);
                       
          assert RAM(1) = "11111110" report "FAIL high bits" severity failure;
          assert RAM(0) = "00000001" report "FAIL low bits" severity failure;
          
        --test #55
          wait for 100 ns;
          wait for c_CLOCK_PERIOD;
          tb_rst <= '1';
          wait for c_CLOCK_PERIOD;
          tb_rst <= '0';
          wait for c_CLOCK_PERIOD;
          tb_start <= '1';
          wait for c_CLOCK_PERIOD;
          tb_start <= '0';
          wait until tb_done = '1';
          wait until tb_done = '0';
          wait until rising_edge(tb_clk);
  
          assert RAM(1) = "11111110" report "FAIL high bits" severity failure;
          assert RAM(0) = "00000001" report "FAIL low bits" severity failure;   
          
        --test #56
            wait for 100 ns;
            wait for c_CLOCK_PERIOD;
            tb_rst <= '1';
            wait for c_CLOCK_PERIOD;
            tb_rst <= '0';
            wait for c_CLOCK_PERIOD;
            tb_start <= '1';
            wait for c_CLOCK_PERIOD;
            tb_start <= '0';
            wait until tb_done = '1';
            wait until tb_done = '0';
            wait until rising_edge(tb_clk);
    
            assert RAM(1) = "11111110" report "FAIL high bits" severity failure;
            assert RAM(0) = "00000001" report "FAIL low bits" severity failure; 
            
        --test #57
              wait for 100 ns;
              wait for c_CLOCK_PERIOD;
              tb_rst <= '1';
              wait for c_CLOCK_PERIOD;
              tb_rst <= '0';
              wait for c_CLOCK_PERIOD;
              tb_start <= '1';
              wait for c_CLOCK_PERIOD;
              tb_start <= '0';
              wait until tb_done = '1';
              wait until tb_done = '0';
              wait until rising_edge(tb_clk);
      
              assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
              assert RAM(0) = "00010000" report "FAIL low bits" severity failure;  
              
        --test #58
                wait for 100 ns;
                wait for c_CLOCK_PERIOD;
                tb_rst <= '1';
                wait for c_CLOCK_PERIOD;
                tb_rst <= '0';
                wait for c_CLOCK_PERIOD;
                tb_start <= '1';
                wait for c_CLOCK_PERIOD;
                tb_start <= '0';
                wait until tb_done = '1';
                wait until tb_done = '0';
                wait until rising_edge(tb_clk);
        
                assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
                assert RAM(0) = "00001001" report "FAIL low bits" severity failure;
                
        --test #59
                wait for 100 ns;
                wait for c_CLOCK_PERIOD;
                tb_rst <= '1';
                wait for c_CLOCK_PERIOD;
                tb_rst <= '0';
                wait for c_CLOCK_PERIOD;
                tb_start <= '1';
                wait for c_CLOCK_PERIOD;
                tb_start <= '0';
                wait until tb_done = '1';
                wait until tb_done = '0';
                wait until rising_edge(tb_clk);
        
                assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
                assert RAM(0) = "00000110" report "FAIL low bits" severity failure;
                
        --test #60
            wait for 100 ns;
            wait for c_CLOCK_PERIOD;
            tb_rst <= '1';
            wait for c_CLOCK_PERIOD;
            tb_rst <= '0';
            wait for c_CLOCK_PERIOD;
            tb_start <= '1';
            wait for c_CLOCK_PERIOD;
            tb_start <= '0';
            wait until tb_done = '1';
            wait until tb_done = '0';
            wait until rising_edge(tb_clk);
    
            assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
            assert RAM(0) = "00000001" report "FAIL low bits" severity failure;
            
        --test #61
            wait for 100 ns;
            wait for c_CLOCK_PERIOD;
            tb_rst <= '1';
            wait for c_CLOCK_PERIOD;
            tb_rst <= '0';
            wait for c_CLOCK_PERIOD;
            tb_start <= '1';
            wait for c_CLOCK_PERIOD;
            tb_start <= '0';
            wait until tb_done = '1';
            wait until tb_done = '0';
            wait until rising_edge(tb_clk);
    
            assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
            assert RAM(0) = "00010000" report "FAIL low bits" severity failure;
            
        --test #62
                wait for 100 ns;
                wait for c_CLOCK_PERIOD;
                tb_rst <= '1';
                wait for c_CLOCK_PERIOD;
                tb_rst <= '0';
                wait for c_CLOCK_PERIOD;
                tb_start <= '1';
                wait for c_CLOCK_PERIOD;
                tb_start <= '0';
                wait until tb_done = '1';
                wait until tb_done = '0';
                wait until rising_edge(tb_clk);
        
                assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
                assert RAM(0) = "00000000" report "FAIL low bits" severity failure;
                
        --test #63
                wait for 100 ns;
                wait for c_CLOCK_PERIOD;
                tb_rst <= '1';
                wait for c_CLOCK_PERIOD;
                tb_rst <= '0';
                wait for c_CLOCK_PERIOD;
                tb_start <= '1';
                wait for c_CLOCK_PERIOD;
                tb_start <= '0';
                wait until tb_done = '1';
                wait until tb_done = '0';
                wait until rising_edge(tb_clk);
        
                assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
                assert RAM(0) = "00000001" report "FAIL low bits" severity failure;
                
        --test #64
                wait for 100 ns;
                wait for c_CLOCK_PERIOD;
                tb_rst <= '1';
                wait for c_CLOCK_PERIOD;
                tb_rst <= '0';
                wait for c_CLOCK_PERIOD;
                tb_start <= '1';
                wait for c_CLOCK_PERIOD;
                tb_start <= '0';
                wait until tb_done = '1';
                wait until tb_done = '0';
                wait until rising_edge(tb_clk);
        
                assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
                assert RAM(0) = "00001100" report "FAIL low bits" severity failure; 
                    
        --test #65
                wait for 100 ns;
                wait for c_CLOCK_PERIOD;
                tb_rst <= '1';
                wait for c_CLOCK_PERIOD;
                tb_rst <= '0';
                wait for c_CLOCK_PERIOD;
                tb_start <= '1';
                wait for c_CLOCK_PERIOD;
                tb_start <= '0';
                wait until tb_done = '1';
                wait until tb_done = '0';
                wait until rising_edge(tb_clk);
        
                assert RAM(1) = "00000000" report "FAIL high bits" severity failure;
                assert RAM(0) = "00000100" report "FAIL low bits" severity failure;                                                                                                                                      




assert false report "Simulation Ended!, test passed" severity failure;
end process test;

end projecttb;